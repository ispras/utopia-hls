module main(	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:11:5
  input  clock,
         reset,
         n_in_0_0_x,
         n_in_0_1_x,
         n_in_0_2_x,
         n_in_0_3_x,
         n_in_0_4_x,
         n_in_0_5_x,
         n_in_0_6_x,
         n_in_0_7_x,
         n_in_1_0_x,
         n_in_1_1_x,
         n_in_1_2_x,
         n_in_1_3_x,
         n_in_1_4_x,
         n_in_1_5_x,
         n_in_1_6_x,
         n_in_1_7_x,
         n_in_2_0_x,
         n_in_2_1_x,
         n_in_2_2_x,
         n_in_2_3_x,
         n_in_2_4_x,
         n_in_2_5_x,
         n_in_2_6_x,
         n_in_2_7_x,
         n_in_3_0_x,
         n_in_3_1_x,
         n_in_3_2_x,
         n_in_3_3_x,
         n_in_3_4_x,
         n_in_3_5_x,
         n_in_3_6_x,
         n_in_3_7_x,
         n_in_4_0_x,
         n_in_4_1_x,
         n_in_4_2_x,
         n_in_4_3_x,
         n_in_4_4_x,
         n_in_4_5_x,
         n_in_4_6_x,
         n_in_4_7_x,
         n_in_5_0_x,
         n_in_5_1_x,
         n_in_5_2_x,
         n_in_5_3_x,
         n_in_5_4_x,
         n_in_5_5_x,
         n_in_5_6_x,
         n_in_5_7_x,
         n_in_6_0_x,
         n_in_6_1_x,
         n_in_6_2_x,
         n_in_6_3_x,
         n_in_6_4_x,
         n_in_6_5_x,
         n_in_6_6_x,
         n_in_6_7_x,
         n_in_7_0_x,
         n_in_7_1_x,
         n_in_7_2_x,
         n_in_7_3_x,
         n_in_7_4_x,
         n_in_7_5_x,
         n_in_7_6_x,
         n_in_7_7_x,
  output n_out_0_0_x,
         n_out_0_1_x,
         n_out_0_2_x,
         n_out_0_3_x,
         n_out_0_4_x,
         n_out_0_5_x,
         n_out_0_6_x,
         n_out_0_7_x,
         n_out_1_0_x,
         n_out_1_1_x,
         n_out_1_2_x,
         n_out_1_3_x,
         n_out_1_4_x,
         n_out_1_5_x,
         n_out_1_6_x,
         n_out_1_7_x,
         n_out_2_0_x,
         n_out_2_1_x,
         n_out_2_2_x,
         n_out_2_3_x,
         n_out_2_4_x,
         n_out_2_5_x,
         n_out_2_6_x,
         n_out_2_7_x,
         n_out_3_0_x,
         n_out_3_1_x,
         n_out_3_2_x,
         n_out_3_3_x,
         n_out_3_4_x,
         n_out_3_5_x,
         n_out_3_6_x,
         n_out_3_7_x,
         n_out_4_0_x,
         n_out_4_1_x,
         n_out_4_2_x,
         n_out_4_3_x,
         n_out_4_4_x,
         n_out_4_5_x,
         n_out_4_6_x,
         n_out_4_7_x,
         n_out_5_0_x,
         n_out_5_1_x,
         n_out_5_2_x,
         n_out_5_3_x,
         n_out_5_4_x,
         n_out_5_5_x,
         n_out_5_6_x,
         n_out_5_7_x,
         n_out_6_0_x,
         n_out_6_1_x,
         n_out_6_2_x,
         n_out_6_3_x,
         n_out_6_4_x,
         n_out_6_5_x,
         n_out_6_6_x,
         n_out_6_7_x,
         n_out_7_0_x,
         n_out_7_1_x,
         n_out_7_2_x,
         n_out_7_3_x,
         n_out_7_4_x,
         n_out_7_5_x,
         n_out_7_6_x,
         n_out_7_7_x);

  wire _delay_INT16_58_2325_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2343:114
  wire _delay_INT16_19_2324_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2342:114
  wire _delay_INT16_49_2323_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2341:114
  wire _delay_INT16_226_2322_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2340:118
  wire _delay_INT16_6_2321_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2339:110
  wire _delay_INT16_23_2320_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2338:114
  wire _delay_INT16_121_2319_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2337:118
  wire _delay_INT16_234_2318_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2336:118
  wire _delay_INT16_132_2317_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2335:118
  wire _delay_INT16_19_2316_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2334:114
  wire _delay_INT16_34_2315_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2333:114
  wire _delay_INT16_378_2314_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2332:118
  wire _delay_INT16_119_2313_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2331:118
  wire _delay_INT16_10_2312_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2330:114
  wire _delay_INT16_158_2311_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2329:118
  wire _delay_INT16_306_2310_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2328:118
  wire _delay_INT16_14_2309_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2327:114
  wire _delay_INT16_230_2308_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2326:118
  wire _delay_INT16_152_2307_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2325:118
  wire _delay_INT16_142_2306_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2324:118
  wire _delay_INT16_180_2305_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2323:118
  wire _delay_INT16_193_2304_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2322:118
  wire _delay_INT16_104_2303_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2321:118
  wire _delay_INT16_2_2302_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2320:110
  wire _delay_INT16_29_2301_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2319:114
  wire _delay_INT16_61_2300_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2318:114
  wire _delay_INT16_268_2299_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2317:118
  wire _delay_INT16_108_2298_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2316:118
  wire _delay_INT16_106_2297_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2315:118
  wire _delay_INT16_7_2296_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2314:110
  wire _delay_INT16_45_2295_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2313:114
  wire _delay_INT16_1_2294_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2312:110
  wire _delay_INT16_200_2293_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2311:118
  wire _delay_INT16_149_2292_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2310:118
  wire _delay_INT16_24_2291_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2309:114
  wire _delay_INT16_171_2290_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2308:118
  wire _delay_INT16_15_2289_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2307:114
  wire _delay_INT16_93_2288_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2306:114
  wire _delay_INT16_29_2287_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2305:114
  wire _delay_INT16_245_2286_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2304:118
  wire _delay_INT16_100_2285_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2303:118
  wire _delay_INT16_350_2284_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2302:118
  wire _delay_INT16_27_2283_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2301:114
  wire _delay_INT16_147_2282_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2300:118
  wire _delay_INT16_127_2281_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2299:118
  wire _delay_INT16_31_2280_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2298:114
  wire _delay_INT16_42_2279_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2297:114
  wire _delay_INT16_137_2278_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2296:118
  wire _delay_INT16_42_2277_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2295:114
  wire _delay_INT16_65_2276_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2294:114
  wire _delay_INT16_65_2275_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2293:114
  wire _delay_INT16_162_2274_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2292:118
  wire _delay_INT16_162_2273_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2291:118
  wire _delay_INT16_120_2272_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2290:118
  wire _delay_INT16_106_2271_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2289:118
  wire _delay_INT16_89_2270_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2288:114
  wire _delay_INT16_89_2269_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2287:114
  wire _delay_INT16_75_2268_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2286:114
  wire _delay_INT16_20_2267_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2285:114
  wire _delay_INT16_206_2266_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2284:118
  wire _delay_INT16_225_2265_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2283:118
  wire _delay_INT16_162_2264_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2282:118
  wire _delay_INT16_49_2263_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2281:114
  wire _delay_INT16_162_2262_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2280:118
  wire _delay_INT16_206_2261_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2279:118
  wire _delay_INT16_20_2260_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2278:114
  wire _delay_INT16_72_2259_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2277:114
  wire _delay_INT16_80_2258_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2276:114
  wire _delay_INT16_23_2257_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2275:114
  wire _delay_INT16_26_2256_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2274:114
  wire _delay_INT16_97_2255_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2273:114
  wire _delay_INT16_14_2254_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2272:114
  wire _delay_INT16_29_2253_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2271:114
  wire _delay_INT16_109_2252_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2270:118
  wire _delay_INT16_6_2251_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2269:110
  wire _delay_INT16_89_2250_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2268:114
  wire _delay_INT16_61_2249_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2267:114
  wire _delay_INT16_83_2248_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2266:114
  wire _delay_INT16_61_2247_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2265:114
  wire _delay_INT16_10_2246_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2264:114
  wire _delay_INT16_139_2245_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2263:118
  wire _delay_INT16_61_2244_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2262:114
  wire _delay_INT16_85_2243_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2261:114
  wire _delay_INT16_85_2242_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2260:114
  wire _delay_INT16_126_2241_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2259:118
  wire _delay_INT16_126_2240_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2258:118
  wire _delay_INT16_85_2239_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2257:114
  wire _delay_INT16_85_2238_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2256:114
  wire _delay_INT16_153_2237_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2255:118
  wire _delay_INT16_153_2236_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2254:118
  wire _delay_INT16_70_2235_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2253:114
  wire _delay_INT16_48_2234_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2252:114
  wire _delay_INT16_48_2233_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2251:114
  wire _delay_INT16_115_2232_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2250:118
  wire _delay_INT16_64_2231_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2249:114
  wire _delay_INT16_100_2230_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2248:118
  wire _delay_INT16_18_2229_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2247:114
  wire _delay_INT16_268_2228_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2246:118
  wire _delay_INT16_303_2227_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2245:118
  wire _delay_INT16_70_2226_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2244:114
  wire _delay_INT16_187_2225_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2243:118
  wire _delay_INT16_235_2224_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2242:118
  wire _delay_INT16_109_2223_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2241:118
  wire _delay_INT16_303_2222_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2240:118
  wire _delay_INT16_268_2221_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2239:118
  wire _delay_INT16_378_2220_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2238:118
  wire _delay_INT16_18_2219_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2237:114
  wire _delay_INT16_180_2218_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2236:118
  wire _delay_INT16_58_2217_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2235:114
  wire _delay_INT16_114_2216_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2234:118
  wire _delay_INT16_36_2215_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2233:114
  wire _delay_INT16_10_2214_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2232:114
  wire _delay_INT16_149_2213_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2231:118
  wire _delay_INT16_289_2212_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2230:118
  wire _delay_INT16_161_2211_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2229:118
  wire _delay_INT16_117_2210_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2228:118
  wire _delay_INT16_217_2209_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2227:118
  wire _delay_INT16_117_2208_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2226:118
  wire _delay_INT16_109_2207_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2225:118
  wire _delay_INT16_106_2206_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2224:118
  wire _delay_INT16_78_2205_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2223:114
  wire _delay_INT16_71_2204_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2222:114
  wire _delay_INT16_74_2203_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2221:114
  wire _delay_INT16_188_2202_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2220:118
  wire _delay_INT16_61_2201_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2219:114
  wire _delay_INT16_34_2200_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2218:114
  wire _delay_INT16_34_2199_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2217:114
  wire _delay_INT16_143_2198_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2216:118
  wire _delay_INT16_143_2197_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2215:118
  wire _delay_INT16_132_2196_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2214:118
  wire _delay_INT16_27_2195_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2213:114
  wire _delay_INT16_180_2194_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2212:118
  wire _delay_INT16_186_2193_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2211:118
  wire _delay_INT16_27_2192_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2210:114
  wire _delay_INT16_72_2191_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2209:114
  wire _delay_INT16_63_2190_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2208:114
  wire _delay_INT16_161_2189_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2207:118
  wire _delay_INT16_72_2188_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2206:114
  wire _delay_INT16_184_2187_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2205:118
  wire _delay_INT16_143_2186_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2204:118
  wire _delay_INT16_184_2185_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2203:118
  wire _delay_INT16_191_2184_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2202:118
  wire _delay_INT16_302_2183_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2201:118
  wire _delay_INT16_10_2182_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2200:114
  wire _delay_INT16_302_2181_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2199:118
  wire _delay_INT16_39_2180_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2198:114
  wire _delay_INT16_191_2179_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2197:118
  wire _delay_INT16_139_2178_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2196:118
  wire _delay_INT16_225_2177_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2195:118
  wire _delay_INT16_143_2176_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2194:118
  wire _delay_INT16_74_2175_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2193:114
  wire _delay_INT16_184_2174_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2192:118
  wire _delay_INT16_16_2173_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2191:114
  wire _delay_INT16_93_2172_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2190:114
  wire _delay_INT16_104_2171_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2189:118
  wire _delay_INT16_40_2170_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2188:114
  wire _delay_INT16_64_2169_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2187:114
  wire _delay_INT16_53_2168_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2186:114
  wire _delay_INT16_60_2167_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2185:114
  wire _delay_INT16_11_2166_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2184:114
  wire _delay_INT16_80_2165_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2183:114
  wire _delay_INT16_206_2164_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2182:118
  wire _delay_INT16_96_2163_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2181:114
  wire _delay_INT16_11_2162_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2180:114
  wire _delay_INT16_11_2161_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2179:114
  wire _delay_INT16_49_2160_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2178:114
  wire _delay_INT16_49_2159_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2177:114
  wire _delay_INT16_119_2158_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2176:118
  wire _delay_INT16_40_2157_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2175:114
  wire _delay_INT16_51_2156_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2174:114
  wire _delay_INT16_125_2155_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2173:118
  wire _delay_INT16_125_2154_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2172:118
  wire _delay_INT16_127_2153_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2171:118
  wire _delay_INT16_157_2152_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2170:118
  wire _delay_INT16_477_2151_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2169:118
  wire _delay_INT16_31_2150_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2168:114
  wire _delay_INT16_152_2149_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2167:118
  wire _delay_INT16_157_2148_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2166:118
  wire _delay_INT16_127_2147_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2165:118
  wire _delay_INT16_48_2146_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2164:114
  wire _delay_INT16_248_2145_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2163:118
  wire _delay_INT16_57_2144_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2162:114
  wire _delay_INT16_60_2143_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2161:114
  wire _delay_INT16_339_2142_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2160:118
  wire _delay_INT16_28_2141_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2159:114
  wire _delay_INT16_24_2140_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2158:114
  wire _delay_INT16_131_2139_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2157:118
  wire _delay_INT16_82_2138_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2156:114
  wire _delay_INT16_26_2137_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2155:114
  wire _delay_INT16_184_2136_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2154:118
  wire _delay_INT16_185_2135_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2153:118
  wire _delay_INT16_145_2134_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2152:118
  wire _delay_INT16_68_2133_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2151:114
  wire _delay_INT16_79_2132_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2150:114
  wire _delay_INT16_79_2131_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2149:114
  wire _delay_INT16_95_2130_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2148:114
  wire _delay_INT16_95_2129_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2147:114
  wire _delay_INT16_229_2128_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2146:118
  wire _delay_INT16_117_2127_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2145:118
  wire _delay_INT16_229_2126_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2144:118
  wire _delay_INT16_166_2125_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2143:118
  wire _delay_INT16_166_2124_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2142:118
  wire _delay_INT16_370_2123_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2141:118
  wire _delay_INT16_114_2122_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2140:118
  wire _delay_INT16_66_2121_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2139:114
  wire _delay_INT16_114_2120_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2138:118
  wire _delay_INT16_83_2119_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2137:114
  wire _delay_INT16_248_2118_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2136:118
  wire _delay_INT16_350_2117_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2135:118
  wire _delay_INT16_141_2116_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2134:118
  wire _delay_INT16_222_2115_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2133:118
  wire _delay_INT16_248_2114_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2132:118
  wire _delay_INT16_83_2113_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2131:114
  wire _delay_INT16_68_2112_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2130:114
  wire _delay_INT16_73_2111_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2129:114
  wire _delay_INT16_87_2110_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2128:114
  wire _delay_INT16_10_2109_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2127:114
  wire _delay_INT16_13_2108_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2126:114
  wire _delay_INT16_121_2107_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2125:118
  wire _delay_INT16_10_2106_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2124:114
  wire _delay_INT16_43_2105_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2123:114
  wire _delay_INT16_87_2104_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2122:114
  wire _delay_INT16_8_2103_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2121:110
  wire _delay_INT16_8_2102_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2120:110
  wire _delay_INT16_31_2101_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2119:114
  wire _delay_INT16_226_2100_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2118:118
  wire _delay_INT16_224_2099_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2117:118
  wire _delay_INT16_5_2098_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2116:110
  wire _delay_INT16_24_2097_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2115:114
  wire _delay_INT16_5_2096_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2114:110
  wire _delay_INT16_61_2095_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2113:114
  wire _delay_INT16_61_2094_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2112:114
  wire _delay_INT16_33_2093_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2111:114
  wire _delay_INT16_115_2092_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2110:118
  wire _delay_INT16_78_2091_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2109:114
  wire _delay_INT16_141_2090_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2108:118
  wire _delay_INT16_63_2089_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2107:114
  wire _delay_INT16_142_2088_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2106:118
  wire _delay_INT16_134_2087_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2105:118
  wire _delay_INT16_134_2086_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2104:118
  wire _delay_INT16_134_2085_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2103:118
  wire _delay_INT16_134_2084_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2102:118
  wire _delay_INT16_131_2083_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2101:118
  wire _delay_INT16_24_2082_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2100:114
  wire _delay_INT16_2_2081_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2099:110
  wire _delay_INT16_1_2080_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2098:110
  wire _delay_INT16_47_2079_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2097:114
  wire _delay_INT16_173_2078_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2096:118
  wire _delay_INT16_3_2077_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2095:110
  wire _delay_INT16_39_2076_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2094:114
  wire _delay_INT16_17_2075_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2093:114
  wire _delay_INT16_11_2074_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2092:114
  wire _delay_INT16_99_2073_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2091:114
  wire _delay_INT16_24_2072_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2090:114
  wire _delay_INT16_24_2071_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2089:114
  wire _delay_INT16_17_2070_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2088:114
  wire _delay_INT16_17_2069_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2087:114
  wire _delay_INT16_15_2068_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2086:114
  wire _delay_INT16_15_2067_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2085:114
  wire _delay_INT16_14_2066_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2084:114
  wire _delay_INT16_14_2065_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2083:114
  wire _delay_INT16_68_2064_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2082:114
  wire _delay_INT16_120_2063_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2081:118
  wire _delay_INT16_396_2062_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2080:118
  wire _delay_INT16_142_2061_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2079:118
  wire _delay_INT16_142_2060_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2078:118
  wire _delay_INT16_339_2059_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2077:118
  wire _delay_INT16_2_2058_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2076:110
  wire _delay_INT16_396_2057_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2075:118
  wire _delay_INT16_50_2056_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2074:114
  wire _delay_INT16_19_2055_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2073:114
  wire _delay_INT16_106_2054_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2072:118
  wire _delay_INT16_34_2053_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2071:114
  wire _delay_INT16_62_2052_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2070:114
  wire _delay_INT16_187_2051_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2069:118
  wire _delay_INT16_111_2050_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2068:118
  wire _delay_INT16_1_2049_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2067:110
  wire _delay_INT16_29_2048_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2066:114
  wire _delay_INT16_182_2047_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2065:118
  wire _delay_INT16_147_2046_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2064:118
  wire _delay_INT16_55_2045_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2063:114
  wire _delay_INT16_48_2044_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2062:114
  wire _delay_INT16_121_2043_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2061:118
  wire _delay_INT16_133_2042_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2060:118
  wire _delay_INT16_13_2041_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2059:114
  wire _delay_INT16_100_2040_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2058:118
  wire _delay_INT16_33_2039_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2057:114
  wire _delay_INT16_35_2038_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2056:114
  wire _delay_INT16_35_2037_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2055:114
  wire _delay_INT16_6_2036_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2054:110
  wire _delay_INT16_19_2035_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2053:114
  wire _delay_INT16_288_2034_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2052:118
  wire _delay_INT16_13_2033_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2051:114
  wire _delay_INT16_13_2032_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2050:114
  wire _delay_INT16_45_2031_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2049:114
  wire _delay_INT16_338_2030_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2048:118
  wire _delay_INT16_255_2029_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2047:118
  wire _delay_INT16_122_2028_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2046:118
  wire _delay_INT16_122_2027_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2045:118
  wire _delay_INT16_255_2026_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2044:118
  wire _delay_INT16_38_2025_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2043:114
  wire _delay_INT16_338_2024_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2042:118
  wire _delay_INT16_45_2023_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2041:114
  wire _delay_INT16_68_2022_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2040:114
  wire _delay_INT16_156_2021_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2039:118
  wire _delay_INT16_64_2020_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2038:114
  wire _delay_INT16_7_2019_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2037:110
  wire _delay_INT16_5_2018_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2036:110
  wire _delay_INT16_298_2017_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2035:118
  wire _delay_INT16_181_2016_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2034:118
  wire _delay_INT16_145_2015_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2033:118
  wire _delay_INT16_242_2014_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2032:118
  wire _delay_INT16_338_2013_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2031:118
  wire _delay_INT16_242_2012_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2030:118
  wire _delay_INT16_127_2011_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2029:118
  wire _delay_INT16_90_2010_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2028:114
  wire _delay_INT16_296_2009_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2027:118
  wire _delay_INT16_81_2008_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2026:114
  wire _delay_INT16_212_2007_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2025:118
  wire _delay_INT16_212_2006_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2024:118
  wire _delay_INT16_21_2005_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2023:114
  wire _delay_INT16_94_2004_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2022:114
  wire _delay_INT16_16_2003_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2021:114
  wire _delay_INT16_94_2002_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2020:114
  wire _delay_INT16_139_2001_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2019:118
  wire _delay_INT16_139_2000_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2018:118
  wire _delay_INT16_23_1999_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2017:114
  wire _delay_INT16_23_1998_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2016:114
  wire _delay_INT16_89_1997_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2015:114
  wire _delay_INT16_89_1996_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2014:114
  wire _delay_INT16_94_1995_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2013:114
  wire _delay_INT16_487_1994_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2012:118
  wire _delay_INT16_34_1993_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2011:114
  wire _delay_INT16_477_1992_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2010:118
  wire _delay_INT16_487_1991_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2009:118
  wire _delay_INT16_94_1990_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2008:114
  wire _delay_INT16_213_1989_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2007:118
  wire _delay_INT16_129_1988_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2006:118
  wire _delay_INT16_262_1987_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2005:118
  wire _delay_INT16_90_1986_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2004:114
  wire _delay_INT16_88_1985_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2003:114
  wire _delay_INT16_259_1984_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2002:118
  wire _delay_INT16_191_1983_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2001:118
  wire _delay_INT16_102_1982_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2000:118
  wire _delay_INT16_131_1981_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1999:118
  wire _delay_INT16_295_1980_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1998:118
  wire _delay_INT16_131_1979_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1997:118
  wire _delay_INT16_397_1978_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1996:118
  wire _delay_INT16_109_1977_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1995:118
  wire _delay_INT16_64_1976_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1994:114
  wire _delay_INT16_10_1975_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1993:114
  wire _delay_INT16_10_1974_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1992:114
  wire _delay_INT16_27_1973_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1991:114
  wire _delay_INT16_27_1972_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1990:114
  wire _delay_INT16_128_1971_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1989:118
  wire _delay_INT16_45_1970_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1988:114
  wire _delay_INT16_45_1969_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1987:114
  wire _delay_INT16_2_1968_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1986:110
  wire _delay_INT16_17_1967_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1985:114
  wire _delay_INT16_1_1966_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1984:110
  wire _delay_INT16_190_1965_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1983:118
  wire _delay_INT16_73_1964_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1982:114
  wire _delay_INT16_19_1963_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1981:114
  wire _delay_INT16_190_1962_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1980:118
  wire _delay_INT16_1_1961_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1979:110
  wire _delay_INT16_2_1960_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1978:110
  wire _delay_INT16_34_1959_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1977:114
  wire _delay_INT16_112_1958_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1976:118
  wire _delay_INT16_68_1957_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1975:114
  wire _delay_INT16_131_1956_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1974:118
  wire _delay_INT16_213_1955_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1973:118
  wire _delay_INT16_66_1954_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1972:114
  wire _delay_INT16_168_1953_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1971:118
  wire _delay_INT16_64_1952_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1970:114
  wire _delay_INT16_75_1951_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1969:114
  wire _delay_INT16_66_1950_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1968:114
  wire _delay_INT16_126_1949_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1967:118
  wire _delay_INT16_1_1948_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1966:110
  wire _delay_INT16_378_1947_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1965:118
  wire _delay_INT16_90_1946_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1964:114
  wire _delay_INT16_122_1945_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1963:118
  wire _delay_INT16_121_1944_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1962:118
  wire _delay_INT16_110_1943_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1961:118
  wire _delay_INT16_145_1942_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1960:118
  wire _delay_INT16_110_1941_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1959:118
  wire _delay_INT16_121_1940_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1958:118
  wire _delay_INT16_122_1939_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1957:118
  wire _delay_INT16_55_1938_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1956:114
  wire _delay_INT16_65_1937_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1955:114
  wire _delay_INT16_178_1936_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1954:118
  wire _delay_INT16_56_1935_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1953:114
  wire _delay_INT16_211_1934_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1952:118
  wire _delay_INT16_176_1933_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1951:118
  wire _delay_INT16_114_1932_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1950:118
  wire _delay_INT16_114_1931_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1949:118
  wire _delay_INT16_1_1930_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1948:110
  wire _delay_INT16_1_1929_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1947:110
  wire _delay_INT16_231_1928_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1946:118
  wire _delay_INT16_59_1927_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1945:114
  wire _delay_INT16_59_1926_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1944:114
  wire _delay_INT16_90_1925_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1943:114
  wire _delay_INT16_90_1924_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1942:114
  wire _delay_INT16_7_1923_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1941:110
  wire _delay_INT16_140_1922_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1940:118
  wire _delay_INT16_106_1921_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1939:118
  wire _delay_INT16_140_1920_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1938:118
  wire _delay_INT16_125_1919_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1937:118
  wire _delay_INT16_125_1918_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1936:118
  wire _delay_INT16_27_1917_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1935:114
  wire _delay_INT16_99_1916_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1934:114
  wire _delay_INT16_351_1915_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1933:118
  wire _delay_INT16_1_1914_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1932:110
  wire _delay_INT16_1_1913_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1931:110
  wire _delay_INT16_222_1912_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1930:118
  wire _delay_INT16_351_1911_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1929:118
  wire _delay_INT16_207_1910_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1928:118
  wire _delay_INT16_159_1909_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1927:118
  wire _delay_INT16_131_1908_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1926:118
  wire _delay_INT16_165_1907_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1925:118
  wire _delay_INT16_165_1906_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1924:118
  wire _delay_INT16_21_1905_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1923:114
  wire _delay_INT16_17_1904_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1922:114
  wire _delay_INT16_38_1903_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1921:114
  wire _delay_INT16_334_1902_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1920:118
  wire _delay_INT16_2_1901_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1919:110
  wire _delay_INT16_334_1900_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1918:118
  wire _delay_INT16_26_1899_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1917:114
  wire _delay_INT16_6_1898_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1916:110
  wire _delay_INT16_14_1897_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1915:114
  wire _delay_INT16_230_1896_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1914:118
  wire _delay_INT16_130_1895_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1913:118
  wire _delay_INT16_121_1894_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1912:118
  wire _delay_INT16_81_1893_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1911:114
  wire _delay_INT16_126_1892_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1910:118
  wire _delay_INT16_378_1891_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1909:118
  wire _delay_INT16_186_1890_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1908:118
  wire _delay_INT16_57_1889_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1907:114
  wire _delay_INT16_57_1888_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1906:114
  wire _delay_INT16_288_1887_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1905:118
  wire _delay_INT16_180_1886_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1904:118
  wire _delay_INT16_11_1885_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1903:114
  wire _delay_INT16_55_1884_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1902:114
  wire _delay_INT16_75_1883_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1901:114
  wire _delay_INT16_5_1882_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1900:110
  wire _delay_INT16_12_1881_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1899:114
  wire _delay_INT16_115_1880_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1898:118
  wire _delay_INT16_81_1879_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1897:114
  wire _delay_INT16_83_1878_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1896:114
  wire _delay_INT16_2_1877_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1895:110
  wire _delay_INT16_128_1876_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1894:118
  wire _delay_INT16_29_1875_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1893:114
  wire _delay_INT16_29_1874_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1892:114
  wire _delay_INT16_126_1873_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1891:118
  wire _delay_INT16_106_1872_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1890:118
  wire _delay_INT16_96_1871_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1889:114
  wire _delay_INT16_136_1870_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1888:118
  wire _delay_INT16_78_1869_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1887:114
  wire _delay_INT16_129_1868_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1886:118
  wire _delay_INT16_86_1867_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1885:114
  wire _delay_INT16_136_1866_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1884:118
  wire _delay_INT16_29_1865_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1883:114
  wire _delay_INT16_1_1864_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1882:110
  wire _delay_INT16_161_1863_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1881:118
  wire _delay_INT16_106_1862_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1880:118
  wire _delay_INT16_106_1861_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1879:118
  wire _delay_INT16_51_1860_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1878:114
  wire _delay_INT16_23_1859_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1877:114
  wire _delay_INT16_23_1858_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1876:114
  wire _delay_INT16_397_1857_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1875:118
  wire _delay_INT16_295_1856_out;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1874:118
  wire _col_7_n_val_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1872:87
  wire _col_7_n_tmp_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1871:105
  wire _col_7_n_val_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1869:87
  wire _col_7_n_tmp_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1868:105
  wire _col_7_n_val_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1866:87
  wire _col_7_n_tmp_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1865:105
  wire _col_7_n_val_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1863:87
  wire _col_7_n_tmp_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1862:105
  wire _col_7_n_val_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1860:87
  wire _col_7_n_tmp_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1859:105
  wire _col_7_n_val_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1857:87
  wire _col_7_n_tmp_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1856:105
  wire _col_7_n_val_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1854:87
  wire _col_7_n_tmp_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1853:105
  wire _col_7_n_val_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1851:87
  wire _col_7_n_tmp_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1850:105
  wire _col_7_d_x4_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1849:100
  wire _col_7_d_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1849:100
  wire _col_7_n_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1848:83
  wire _col_7_n_w4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1847:100
  wire _col_7_n_v4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1846:100
  wire _col_7_n_u4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1845:100
  wire _col_7_d_x2_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1844:100
  wire _col_7_d_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1844:100
  wire _col_7_n_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1843:83
  wire _col_7_n_w2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1842:100
  wire _col_7_n_v2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1841:100
  wire _col_7_n_u2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1840:100
  wire _col_7_d_x0_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1839:100
  wire _col_7_d_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1839:100
  wire _col_7_n_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1838:100
  wire _col_7_d_x3_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1837:100
  wire _col_7_d_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1837:100
  wire _col_7_n_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1836:100
  wire _col_7_d_x8_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1835:100
  wire _col_7_d_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1835:100
  wire _col_7_n_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1834:100
  wire _col_7_d_x7_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1833:100
  wire _col_7_d_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1833:100
  wire _col_7_n_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1832:100
  wire _col_7_d_x5_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1831:100
  wire _col_7_d_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1831:100
  wire _col_7_n_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1830:100
  wire _col_7_d_x6_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1829:100
  wire _col_7_d_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1829:100
  wire _col_7_n_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1828:100
  wire _col_7_d_x4_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1827:100
  wire _col_7_d_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1827:100
  wire _col_7_n_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1826:100
  wire _col_7_d_x1_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1825:100
  wire _col_7_d_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1825:100
  wire _col_7_n_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1824:100
  wire _col_7_d_x3_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1823:100
  wire _col_7_d_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1823:100
  wire _col_7_n_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1822:83
  wire _col_7_n_v3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1821:100
  wire _col_7_n_u3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1820:100
  wire _col_7_d_x2_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1819:100
  wire _col_7_d_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1819:100
  wire _col_7_n_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1818:83
  wire _col_7_n_v2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1817:100
  wire _col_7_n_u2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1816:100
  wire _col_7_d_x1_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1815:100
  wire _col_7_d_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1815:100
  wire _col_7_n_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1814:100
  wire _col_7_n_v1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1813:100
  wire _col_7_n_u1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1812:100
  wire _col_7_d_x0_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1811:100
  wire _col_7_d_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1811:100
  wire _col_7_n_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1810:100
  wire _col_7_d_x8_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1809:100
  wire _col_7_d_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1809:100
  wire _col_7_n_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1808:100
  wire _col_7_d_x7_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1807:100
  wire _col_7_d_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1807:100
  wire _col_7_n_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1806:83
  wire _col_7_n_v7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1805:100
  wire _col_7_n_u7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1804:100
  wire _col_7_d_x6_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1803:100
  wire _col_7_d_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1803:100
  wire _col_7_n_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1802:83
  wire _col_7_n_v6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1801:100
  wire _col_7_n_u6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1800:100
  wire _col_7_d_x8_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1799:100
  wire _col_7_d_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1799:100
  wire _col_7_n_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1798:100
  wire _col_7_n_v8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1797:100
  wire _col_7_n_u8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1796:100
  wire _col_7_d_x5_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1795:100
  wire _col_7_d_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1795:100
  wire _col_7_n_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1794:83
  wire _col_7_n_v5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1793:100
  wire _col_7_n_u5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1792:100
  wire _col_7_d_x4_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1791:100
  wire _col_7_d_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1791:100
  wire _col_7_n_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1790:83
  wire _col_7_n_v4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1789:100
  wire _col_7_n_u4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1788:100
  wire _col_7_d_x8_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1787:100
  wire _col_7_d_x8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1787:100
  wire _col_7_n_x8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1786:100
  wire _col_7_n_v8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1785:100
  wire _col_7_n_u8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1784:100
  wire _col_7_d_x7_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1783:100
  wire _col_7_d_x7_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1783:100
  wire _col_7_d_x6_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1782:100
  wire _col_7_d_x6_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1782:100
  wire _col_7_d_x5_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1781:100
  wire _col_7_d_x5_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1781:100
  wire _col_7_d_x4_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1780:100
  wire _col_7_d_x4_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1780:100
  wire _col_7_d_x3_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1779:100
  wire _col_7_d_x3_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1779:100
  wire _col_7_d_x2_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1778:100
  wire _col_7_d_x2_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1778:100
  wire _col_7_d_x1_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1777:100
  wire _col_7_d_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1777:100
  wire _col_7_d_x0_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1776:100
  wire _col_7_d_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1776:100
  wire _col_7_n_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1775:100
  wire _col_7_n_t0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1774:83
  wire _col_7_n_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1773:83
  wire _col_7_n_w2_add_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1772:85
  wire _col_7_n_w2_sub_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1771:85
  wire _col_7_n_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1770:64
  wire _col_7_n_w3_add_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1769:85
  wire _col_7_n_w3_sub_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1768:85
  wire _col_7_n_w3_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1767:64
  wire _col_7_n_w1_add_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1766:85
  wire _col_7_n_w1_sub_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1765:85
  wire _col_7_n_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1764:64
  wire _col_7_n_c8192_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1763:73
  wire _col_7_n_c181_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1762:76
  wire _col_7_n_c181_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1761:76
  wire _col_7_n_c128_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1760:76
  wire _col_7_n_c128_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1759:76
  wire _col_7_n_c4_2_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1758:70
  wire _col_7_n_c4_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1757:70
  wire _col_7_n_c4_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1756:70
  wire _col_6_n_val_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1754:87
  wire _col_6_n_tmp_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1753:105
  wire _col_6_n_val_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1751:87
  wire _col_6_n_tmp_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1750:105
  wire _col_6_n_val_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1748:87
  wire _col_6_n_tmp_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1747:105
  wire _col_6_n_val_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1745:87
  wire _col_6_n_tmp_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1744:105
  wire _col_6_n_val_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1742:87
  wire _col_6_n_tmp_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1741:105
  wire _col_6_n_val_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1739:87
  wire _col_6_n_tmp_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1738:105
  wire _col_6_n_val_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1736:87
  wire _col_6_n_tmp_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1735:105
  wire _col_6_n_val_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1733:87
  wire _col_6_n_tmp_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1732:105
  wire _col_6_d_x4_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1731:100
  wire _col_6_d_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1731:100
  wire _col_6_n_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1730:83
  wire _col_6_n_w4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1729:100
  wire _col_6_n_v4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1728:100
  wire _col_6_n_u4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1727:100
  wire _col_6_d_x2_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1726:100
  wire _col_6_d_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1726:100
  wire _col_6_n_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1725:83
  wire _col_6_n_w2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1724:100
  wire _col_6_n_v2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1723:100
  wire _col_6_n_u2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1722:100
  wire _col_6_d_x0_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1721:100
  wire _col_6_d_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1721:100
  wire _col_6_n_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1720:100
  wire _col_6_d_x3_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1719:100
  wire _col_6_d_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1719:100
  wire _col_6_n_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1718:100
  wire _col_6_d_x8_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1717:100
  wire _col_6_d_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1717:100
  wire _col_6_n_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1716:100
  wire _col_6_d_x7_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1715:100
  wire _col_6_d_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1715:100
  wire _col_6_n_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1714:100
  wire _col_6_d_x5_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1713:100
  wire _col_6_d_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1713:100
  wire _col_6_n_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1712:100
  wire _col_6_d_x6_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1711:100
  wire _col_6_d_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1711:100
  wire _col_6_n_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1710:100
  wire _col_6_d_x4_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1709:100
  wire _col_6_d_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1709:100
  wire _col_6_n_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1708:100
  wire _col_6_d_x1_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1707:100
  wire _col_6_d_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1707:100
  wire _col_6_n_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1706:100
  wire _col_6_d_x3_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1705:100
  wire _col_6_d_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1705:100
  wire _col_6_n_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1704:83
  wire _col_6_n_v3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1703:100
  wire _col_6_n_u3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1702:100
  wire _col_6_d_x2_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1701:100
  wire _col_6_d_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1701:100
  wire _col_6_n_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1700:83
  wire _col_6_n_v2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1699:100
  wire _col_6_n_u2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1698:100
  wire _col_6_d_x1_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1697:100
  wire _col_6_d_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1697:100
  wire _col_6_n_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1696:100
  wire _col_6_n_v1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1695:100
  wire _col_6_n_u1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1694:100
  wire _col_6_d_x0_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1693:100
  wire _col_6_d_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1693:100
  wire _col_6_n_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1692:100
  wire _col_6_d_x8_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1691:100
  wire _col_6_d_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1691:100
  wire _col_6_n_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1690:100
  wire _col_6_d_x7_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1689:100
  wire _col_6_d_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1689:100
  wire _col_6_n_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1688:83
  wire _col_6_n_v7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1687:100
  wire _col_6_n_u7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1686:100
  wire _col_6_d_x6_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1685:100
  wire _col_6_d_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1685:100
  wire _col_6_n_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1684:83
  wire _col_6_n_v6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1683:100
  wire _col_6_n_u6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1682:100
  wire _col_6_d_x8_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1681:100
  wire _col_6_d_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1681:100
  wire _col_6_n_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1680:100
  wire _col_6_n_v8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1679:100
  wire _col_6_n_u8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1678:100
  wire _col_6_d_x5_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1677:100
  wire _col_6_d_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1677:100
  wire _col_6_n_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1676:83
  wire _col_6_n_v5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1675:100
  wire _col_6_n_u5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1674:100
  wire _col_6_d_x4_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1673:100
  wire _col_6_d_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1673:100
  wire _col_6_n_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1672:83
  wire _col_6_n_v4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1671:100
  wire _col_6_n_u4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1670:100
  wire _col_6_d_x8_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1669:100
  wire _col_6_d_x8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1669:100
  wire _col_6_n_x8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1668:100
  wire _col_6_n_v8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1667:100
  wire _col_6_n_u8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1666:100
  wire _col_6_d_x7_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1665:100
  wire _col_6_d_x7_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1665:100
  wire _col_6_d_x6_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1664:100
  wire _col_6_d_x6_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1664:100
  wire _col_6_d_x5_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1663:100
  wire _col_6_d_x5_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1663:100
  wire _col_6_d_x4_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1662:100
  wire _col_6_d_x4_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1662:100
  wire _col_6_d_x3_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1661:100
  wire _col_6_d_x3_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1661:100
  wire _col_6_d_x2_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1660:100
  wire _col_6_d_x2_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1660:100
  wire _col_6_d_x1_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1659:100
  wire _col_6_d_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1659:100
  wire _col_6_d_x0_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1658:100
  wire _col_6_d_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1658:100
  wire _col_6_n_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1657:100
  wire _col_6_n_t0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1656:83
  wire _col_6_n_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1655:83
  wire _col_6_n_w2_add_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1654:85
  wire _col_6_n_w2_sub_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1653:85
  wire _col_6_n_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1652:64
  wire _col_6_n_w3_add_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1651:85
  wire _col_6_n_w3_sub_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1650:85
  wire _col_6_n_w3_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1649:64
  wire _col_6_n_w1_add_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1648:85
  wire _col_6_n_w1_sub_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1647:85
  wire _col_6_n_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1646:64
  wire _col_6_n_c8192_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1645:73
  wire _col_6_n_c181_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1644:76
  wire _col_6_n_c181_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1643:76
  wire _col_6_n_c128_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1642:76
  wire _col_6_n_c128_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1641:76
  wire _col_6_n_c4_2_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1640:70
  wire _col_6_n_c4_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1639:70
  wire _col_6_n_c4_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1638:70
  wire _col_5_n_val_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1636:87
  wire _col_5_n_tmp_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1635:105
  wire _col_5_n_val_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1633:87
  wire _col_5_n_tmp_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1632:105
  wire _col_5_n_val_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1630:87
  wire _col_5_n_tmp_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1629:105
  wire _col_5_n_val_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1627:87
  wire _col_5_n_tmp_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1626:105
  wire _col_5_n_val_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1624:87
  wire _col_5_n_tmp_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1623:105
  wire _col_5_n_val_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1621:87
  wire _col_5_n_tmp_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1620:105
  wire _col_5_n_val_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1618:87
  wire _col_5_n_tmp_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1617:105
  wire _col_5_n_val_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1615:87
  wire _col_5_n_tmp_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1614:105
  wire _col_5_d_x4_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1613:100
  wire _col_5_d_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1613:100
  wire _col_5_n_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1612:83
  wire _col_5_n_w4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1611:100
  wire _col_5_n_v4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1610:100
  wire _col_5_n_u4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1609:100
  wire _col_5_d_x2_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1608:100
  wire _col_5_d_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1608:100
  wire _col_5_n_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1607:83
  wire _col_5_n_w2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1606:100
  wire _col_5_n_v2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1605:100
  wire _col_5_n_u2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1604:100
  wire _col_5_d_x0_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1603:100
  wire _col_5_d_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1603:100
  wire _col_5_n_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1602:100
  wire _col_5_d_x3_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1601:100
  wire _col_5_d_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1601:100
  wire _col_5_n_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1600:100
  wire _col_5_d_x8_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1599:100
  wire _col_5_d_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1599:100
  wire _col_5_n_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1598:100
  wire _col_5_d_x7_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1597:100
  wire _col_5_d_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1597:100
  wire _col_5_n_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1596:100
  wire _col_5_d_x5_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1595:100
  wire _col_5_d_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1595:100
  wire _col_5_n_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1594:100
  wire _col_5_d_x6_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1593:100
  wire _col_5_d_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1593:100
  wire _col_5_n_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1592:100
  wire _col_5_d_x4_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1591:100
  wire _col_5_d_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1591:100
  wire _col_5_n_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1590:100
  wire _col_5_d_x1_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1589:100
  wire _col_5_d_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1589:100
  wire _col_5_n_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1588:100
  wire _col_5_d_x3_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1587:100
  wire _col_5_d_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1587:100
  wire _col_5_n_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1586:83
  wire _col_5_n_v3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1585:100
  wire _col_5_n_u3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1584:100
  wire _col_5_d_x2_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1583:100
  wire _col_5_d_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1583:100
  wire _col_5_n_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1582:83
  wire _col_5_n_v2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1581:100
  wire _col_5_n_u2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1580:100
  wire _col_5_d_x1_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1579:100
  wire _col_5_d_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1579:100
  wire _col_5_n_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1578:100
  wire _col_5_n_v1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1577:100
  wire _col_5_n_u1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1576:100
  wire _col_5_d_x0_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1575:100
  wire _col_5_d_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1575:100
  wire _col_5_n_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1574:100
  wire _col_5_d_x8_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1573:100
  wire _col_5_d_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1573:100
  wire _col_5_n_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1572:100
  wire _col_5_d_x7_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1571:100
  wire _col_5_d_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1571:100
  wire _col_5_n_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1570:83
  wire _col_5_n_v7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1569:100
  wire _col_5_n_u7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1568:100
  wire _col_5_d_x6_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1567:100
  wire _col_5_d_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1567:100
  wire _col_5_n_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1566:83
  wire _col_5_n_v6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1565:100
  wire _col_5_n_u6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1564:100
  wire _col_5_d_x8_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1563:100
  wire _col_5_d_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1563:100
  wire _col_5_n_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1562:100
  wire _col_5_n_v8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1561:100
  wire _col_5_n_u8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1560:100
  wire _col_5_d_x5_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1559:100
  wire _col_5_d_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1559:100
  wire _col_5_n_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1558:83
  wire _col_5_n_v5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1557:100
  wire _col_5_n_u5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1556:100
  wire _col_5_d_x4_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1555:100
  wire _col_5_d_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1555:100
  wire _col_5_n_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1554:83
  wire _col_5_n_v4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1553:100
  wire _col_5_n_u4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1552:100
  wire _col_5_d_x8_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1551:100
  wire _col_5_d_x8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1551:100
  wire _col_5_n_x8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1550:100
  wire _col_5_n_v8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1549:100
  wire _col_5_n_u8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1548:100
  wire _col_5_d_x7_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1547:100
  wire _col_5_d_x7_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1547:100
  wire _col_5_d_x6_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1546:100
  wire _col_5_d_x6_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1546:100
  wire _col_5_d_x5_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1545:100
  wire _col_5_d_x5_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1545:100
  wire _col_5_d_x4_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1544:100
  wire _col_5_d_x4_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1544:100
  wire _col_5_d_x3_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1543:100
  wire _col_5_d_x3_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1543:100
  wire _col_5_d_x2_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1542:100
  wire _col_5_d_x2_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1542:100
  wire _col_5_d_x1_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1541:100
  wire _col_5_d_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1541:100
  wire _col_5_d_x0_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1540:100
  wire _col_5_d_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1540:100
  wire _col_5_n_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1539:100
  wire _col_5_n_t0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1538:83
  wire _col_5_n_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1537:83
  wire _col_5_n_w2_add_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1536:85
  wire _col_5_n_w2_sub_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1535:85
  wire _col_5_n_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1534:64
  wire _col_5_n_w3_add_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1533:85
  wire _col_5_n_w3_sub_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1532:85
  wire _col_5_n_w3_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1531:64
  wire _col_5_n_w1_add_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1530:85
  wire _col_5_n_w1_sub_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1529:85
  wire _col_5_n_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1528:64
  wire _col_5_n_c8192_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1527:73
  wire _col_5_n_c181_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1526:76
  wire _col_5_n_c181_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1525:76
  wire _col_5_n_c128_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1524:76
  wire _col_5_n_c128_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1523:76
  wire _col_5_n_c4_2_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1522:70
  wire _col_5_n_c4_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1521:70
  wire _col_5_n_c4_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1520:70
  wire _col_4_n_val_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1518:87
  wire _col_4_n_tmp_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1517:105
  wire _col_4_n_val_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1515:87
  wire _col_4_n_tmp_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1514:105
  wire _col_4_n_val_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1512:87
  wire _col_4_n_tmp_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1511:105
  wire _col_4_n_val_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1509:87
  wire _col_4_n_tmp_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1508:105
  wire _col_4_n_val_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1506:87
  wire _col_4_n_tmp_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1505:105
  wire _col_4_n_val_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1503:87
  wire _col_4_n_tmp_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1502:105
  wire _col_4_n_val_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1500:87
  wire _col_4_n_tmp_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1499:105
  wire _col_4_n_val_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1497:87
  wire _col_4_n_tmp_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1496:105
  wire _col_4_d_x4_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1495:100
  wire _col_4_d_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1495:100
  wire _col_4_n_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1494:83
  wire _col_4_n_w4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1493:100
  wire _col_4_n_v4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1492:100
  wire _col_4_n_u4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1491:100
  wire _col_4_d_x2_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1490:100
  wire _col_4_d_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1490:100
  wire _col_4_n_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1489:83
  wire _col_4_n_w2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1488:100
  wire _col_4_n_v2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1487:100
  wire _col_4_n_u2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1486:100
  wire _col_4_d_x0_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1485:100
  wire _col_4_d_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1485:100
  wire _col_4_n_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1484:100
  wire _col_4_d_x3_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1483:100
  wire _col_4_d_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1483:100
  wire _col_4_n_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1482:100
  wire _col_4_d_x8_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1481:100
  wire _col_4_d_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1481:100
  wire _col_4_n_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1480:100
  wire _col_4_d_x7_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1479:100
  wire _col_4_d_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1479:100
  wire _col_4_n_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1478:100
  wire _col_4_d_x5_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1477:100
  wire _col_4_d_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1477:100
  wire _col_4_n_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1476:100
  wire _col_4_d_x6_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1475:100
  wire _col_4_d_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1475:100
  wire _col_4_n_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1474:100
  wire _col_4_d_x4_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1473:100
  wire _col_4_d_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1473:100
  wire _col_4_n_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1472:100
  wire _col_4_d_x1_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1471:100
  wire _col_4_d_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1471:100
  wire _col_4_n_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1470:100
  wire _col_4_d_x3_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1469:100
  wire _col_4_d_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1469:100
  wire _col_4_n_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1468:83
  wire _col_4_n_v3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1467:100
  wire _col_4_n_u3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1466:100
  wire _col_4_d_x2_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1465:100
  wire _col_4_d_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1465:100
  wire _col_4_n_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1464:83
  wire _col_4_n_v2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1463:100
  wire _col_4_n_u2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1462:100
  wire _col_4_d_x1_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1461:100
  wire _col_4_d_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1461:100
  wire _col_4_n_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1460:100
  wire _col_4_n_v1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1459:100
  wire _col_4_n_u1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1458:100
  wire _col_4_d_x0_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1457:100
  wire _col_4_d_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1457:100
  wire _col_4_n_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1456:100
  wire _col_4_d_x8_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1455:100
  wire _col_4_d_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1455:100
  wire _col_4_n_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1454:100
  wire _col_4_d_x7_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1453:100
  wire _col_4_d_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1453:100
  wire _col_4_n_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1452:83
  wire _col_4_n_v7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1451:100
  wire _col_4_n_u7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1450:100
  wire _col_4_d_x6_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1449:100
  wire _col_4_d_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1449:100
  wire _col_4_n_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1448:83
  wire _col_4_n_v6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1447:100
  wire _col_4_n_u6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1446:100
  wire _col_4_d_x8_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1445:100
  wire _col_4_d_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1445:100
  wire _col_4_n_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1444:100
  wire _col_4_n_v8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1443:100
  wire _col_4_n_u8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1442:100
  wire _col_4_d_x5_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1441:100
  wire _col_4_d_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1441:100
  wire _col_4_n_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1440:83
  wire _col_4_n_v5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1439:100
  wire _col_4_n_u5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1438:100
  wire _col_4_d_x4_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1437:100
  wire _col_4_d_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1437:100
  wire _col_4_n_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1436:83
  wire _col_4_n_v4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1435:100
  wire _col_4_n_u4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1434:100
  wire _col_4_d_x8_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1433:100
  wire _col_4_d_x8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1433:100
  wire _col_4_n_x8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1432:100
  wire _col_4_n_v8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1431:100
  wire _col_4_n_u8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1430:100
  wire _col_4_d_x7_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1429:100
  wire _col_4_d_x7_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1429:100
  wire _col_4_d_x6_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1428:100
  wire _col_4_d_x6_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1428:100
  wire _col_4_d_x5_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1427:100
  wire _col_4_d_x5_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1427:100
  wire _col_4_d_x4_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1426:100
  wire _col_4_d_x4_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1426:100
  wire _col_4_d_x3_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1425:100
  wire _col_4_d_x3_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1425:100
  wire _col_4_d_x2_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1424:100
  wire _col_4_d_x2_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1424:100
  wire _col_4_d_x1_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1423:100
  wire _col_4_d_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1423:100
  wire _col_4_d_x0_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1422:100
  wire _col_4_d_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1422:100
  wire _col_4_n_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1421:100
  wire _col_4_n_t0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1420:83
  wire _col_4_n_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1419:83
  wire _col_4_n_w2_add_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1418:85
  wire _col_4_n_w2_sub_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1417:85
  wire _col_4_n_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1416:64
  wire _col_4_n_w3_add_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1415:85
  wire _col_4_n_w3_sub_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1414:85
  wire _col_4_n_w3_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1413:64
  wire _col_4_n_w1_add_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1412:85
  wire _col_4_n_w1_sub_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1411:85
  wire _col_4_n_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1410:64
  wire _col_4_n_c8192_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1409:73
  wire _col_4_n_c181_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1408:76
  wire _col_4_n_c181_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1407:76
  wire _col_4_n_c128_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1406:76
  wire _col_4_n_c128_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1405:76
  wire _col_4_n_c4_2_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1404:70
  wire _col_4_n_c4_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1403:70
  wire _col_4_n_c4_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1402:70
  wire _col_3_n_val_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1400:87
  wire _col_3_n_tmp_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1399:105
  wire _col_3_n_val_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1397:87
  wire _col_3_n_tmp_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1396:105
  wire _col_3_n_val_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1394:87
  wire _col_3_n_tmp_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1393:105
  wire _col_3_n_val_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1391:87
  wire _col_3_n_tmp_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1390:105
  wire _col_3_n_val_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1388:87
  wire _col_3_n_tmp_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1387:105
  wire _col_3_n_val_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1385:87
  wire _col_3_n_tmp_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1384:105
  wire _col_3_n_val_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1382:87
  wire _col_3_n_tmp_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1381:105
  wire _col_3_n_val_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1379:87
  wire _col_3_n_tmp_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1378:105
  wire _col_3_d_x4_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1377:100
  wire _col_3_d_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1377:100
  wire _col_3_n_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1376:83
  wire _col_3_n_w4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1375:100
  wire _col_3_n_v4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1374:100
  wire _col_3_n_u4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1373:100
  wire _col_3_d_x2_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1372:100
  wire _col_3_d_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1372:100
  wire _col_3_n_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1371:83
  wire _col_3_n_w2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1370:100
  wire _col_3_n_v2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1369:100
  wire _col_3_n_u2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1368:100
  wire _col_3_d_x0_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1367:100
  wire _col_3_d_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1367:100
  wire _col_3_n_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1366:100
  wire _col_3_d_x3_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1365:100
  wire _col_3_d_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1365:100
  wire _col_3_n_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1364:100
  wire _col_3_d_x8_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1363:100
  wire _col_3_d_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1363:100
  wire _col_3_n_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1362:100
  wire _col_3_d_x7_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1361:100
  wire _col_3_d_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1361:100
  wire _col_3_n_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1360:100
  wire _col_3_d_x5_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1359:100
  wire _col_3_d_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1359:100
  wire _col_3_n_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1358:100
  wire _col_3_d_x6_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1357:100
  wire _col_3_d_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1357:100
  wire _col_3_n_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1356:100
  wire _col_3_d_x4_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1355:100
  wire _col_3_d_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1355:100
  wire _col_3_n_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1354:100
  wire _col_3_d_x1_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1353:100
  wire _col_3_d_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1353:100
  wire _col_3_n_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1352:100
  wire _col_3_d_x3_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1351:100
  wire _col_3_d_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1351:100
  wire _col_3_n_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1350:83
  wire _col_3_n_v3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1349:100
  wire _col_3_n_u3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1348:100
  wire _col_3_d_x2_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1347:100
  wire _col_3_d_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1347:100
  wire _col_3_n_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1346:83
  wire _col_3_n_v2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1345:100
  wire _col_3_n_u2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1344:100
  wire _col_3_d_x1_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1343:100
  wire _col_3_d_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1343:100
  wire _col_3_n_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1342:100
  wire _col_3_n_v1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1341:100
  wire _col_3_n_u1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1340:100
  wire _col_3_d_x0_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1339:100
  wire _col_3_d_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1339:100
  wire _col_3_n_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1338:100
  wire _col_3_d_x8_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1337:100
  wire _col_3_d_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1337:100
  wire _col_3_n_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1336:100
  wire _col_3_d_x7_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1335:100
  wire _col_3_d_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1335:100
  wire _col_3_n_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1334:83
  wire _col_3_n_v7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1333:100
  wire _col_3_n_u7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1332:100
  wire _col_3_d_x6_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1331:100
  wire _col_3_d_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1331:100
  wire _col_3_n_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1330:83
  wire _col_3_n_v6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1329:100
  wire _col_3_n_u6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1328:100
  wire _col_3_d_x8_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1327:100
  wire _col_3_d_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1327:100
  wire _col_3_n_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1326:100
  wire _col_3_n_v8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1325:100
  wire _col_3_n_u8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1324:100
  wire _col_3_d_x5_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1323:100
  wire _col_3_d_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1323:100
  wire _col_3_n_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1322:83
  wire _col_3_n_v5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1321:100
  wire _col_3_n_u5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1320:100
  wire _col_3_d_x4_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1319:100
  wire _col_3_d_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1319:100
  wire _col_3_n_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1318:83
  wire _col_3_n_v4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1317:100
  wire _col_3_n_u4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1316:100
  wire _col_3_d_x8_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1315:100
  wire _col_3_d_x8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1315:100
  wire _col_3_n_x8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1314:100
  wire _col_3_n_v8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1313:100
  wire _col_3_n_u8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1312:100
  wire _col_3_d_x7_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1311:100
  wire _col_3_d_x7_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1311:100
  wire _col_3_d_x6_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1310:100
  wire _col_3_d_x6_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1310:100
  wire _col_3_d_x5_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1309:100
  wire _col_3_d_x5_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1309:100
  wire _col_3_d_x4_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1308:100
  wire _col_3_d_x4_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1308:100
  wire _col_3_d_x3_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1307:100
  wire _col_3_d_x3_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1307:100
  wire _col_3_d_x2_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1306:100
  wire _col_3_d_x2_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1306:100
  wire _col_3_d_x1_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1305:100
  wire _col_3_d_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1305:100
  wire _col_3_d_x0_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1304:100
  wire _col_3_d_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1304:100
  wire _col_3_n_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1303:100
  wire _col_3_n_t0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1302:83
  wire _col_3_n_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1301:83
  wire _col_3_n_w2_add_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1300:85
  wire _col_3_n_w2_sub_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1299:85
  wire _col_3_n_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1298:64
  wire _col_3_n_w3_add_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1297:85
  wire _col_3_n_w3_sub_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1296:85
  wire _col_3_n_w3_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1295:64
  wire _col_3_n_w1_add_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1294:85
  wire _col_3_n_w1_sub_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1293:85
  wire _col_3_n_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1292:64
  wire _col_3_n_c8192_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1291:73
  wire _col_3_n_c181_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1290:76
  wire _col_3_n_c181_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1289:76
  wire _col_3_n_c128_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1288:76
  wire _col_3_n_c128_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1287:76
  wire _col_3_n_c4_2_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1286:70
  wire _col_3_n_c4_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1285:70
  wire _col_3_n_c4_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1284:70
  wire _col_2_n_val_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1282:87
  wire _col_2_n_tmp_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1281:105
  wire _col_2_n_val_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1279:87
  wire _col_2_n_tmp_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1278:105
  wire _col_2_n_val_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1276:87
  wire _col_2_n_tmp_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1275:105
  wire _col_2_n_val_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1273:87
  wire _col_2_n_tmp_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1272:105
  wire _col_2_n_val_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1270:87
  wire _col_2_n_tmp_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1269:105
  wire _col_2_n_val_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1267:87
  wire _col_2_n_tmp_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1266:105
  wire _col_2_n_val_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1264:87
  wire _col_2_n_tmp_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1263:105
  wire _col_2_n_val_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1261:87
  wire _col_2_n_tmp_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1260:105
  wire _col_2_d_x4_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1259:100
  wire _col_2_d_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1259:100
  wire _col_2_n_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1258:83
  wire _col_2_n_w4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1257:100
  wire _col_2_n_v4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1256:100
  wire _col_2_n_u4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1255:100
  wire _col_2_d_x2_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1254:100
  wire _col_2_d_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1254:100
  wire _col_2_n_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1253:83
  wire _col_2_n_w2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1252:100
  wire _col_2_n_v2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1251:100
  wire _col_2_n_u2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1250:100
  wire _col_2_d_x0_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1249:100
  wire _col_2_d_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1249:100
  wire _col_2_n_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1248:100
  wire _col_2_d_x3_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1247:100
  wire _col_2_d_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1247:100
  wire _col_2_n_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1246:100
  wire _col_2_d_x8_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1245:100
  wire _col_2_d_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1245:100
  wire _col_2_n_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1244:100
  wire _col_2_d_x7_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1243:100
  wire _col_2_d_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1243:100
  wire _col_2_n_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1242:100
  wire _col_2_d_x5_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1241:100
  wire _col_2_d_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1241:100
  wire _col_2_n_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1240:100
  wire _col_2_d_x6_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1239:100
  wire _col_2_d_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1239:100
  wire _col_2_n_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1238:100
  wire _col_2_d_x4_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1237:100
  wire _col_2_d_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1237:100
  wire _col_2_n_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1236:100
  wire _col_2_d_x1_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1235:100
  wire _col_2_d_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1235:100
  wire _col_2_n_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1234:100
  wire _col_2_d_x3_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1233:100
  wire _col_2_d_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1233:100
  wire _col_2_n_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1232:83
  wire _col_2_n_v3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1231:100
  wire _col_2_n_u3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1230:100
  wire _col_2_d_x2_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1229:100
  wire _col_2_d_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1229:100
  wire _col_2_n_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1228:83
  wire _col_2_n_v2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1227:100
  wire _col_2_n_u2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1226:100
  wire _col_2_d_x1_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1225:100
  wire _col_2_d_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1225:100
  wire _col_2_n_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1224:100
  wire _col_2_n_v1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1223:100
  wire _col_2_n_u1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1222:100
  wire _col_2_d_x0_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1221:100
  wire _col_2_d_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1221:100
  wire _col_2_n_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1220:100
  wire _col_2_d_x8_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1219:100
  wire _col_2_d_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1219:100
  wire _col_2_n_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1218:100
  wire _col_2_d_x7_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1217:100
  wire _col_2_d_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1217:100
  wire _col_2_n_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1216:83
  wire _col_2_n_v7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1215:100
  wire _col_2_n_u7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1214:100
  wire _col_2_d_x6_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1213:100
  wire _col_2_d_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1213:100
  wire _col_2_n_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1212:83
  wire _col_2_n_v6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1211:100
  wire _col_2_n_u6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1210:100
  wire _col_2_d_x8_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1209:100
  wire _col_2_d_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1209:100
  wire _col_2_n_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1208:100
  wire _col_2_n_v8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1207:100
  wire _col_2_n_u8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1206:100
  wire _col_2_d_x5_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1205:100
  wire _col_2_d_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1205:100
  wire _col_2_n_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1204:83
  wire _col_2_n_v5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1203:100
  wire _col_2_n_u5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1202:100
  wire _col_2_d_x4_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1201:100
  wire _col_2_d_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1201:100
  wire _col_2_n_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1200:83
  wire _col_2_n_v4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1199:100
  wire _col_2_n_u4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1198:100
  wire _col_2_d_x8_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1197:100
  wire _col_2_d_x8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1197:100
  wire _col_2_n_x8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1196:100
  wire _col_2_n_v8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1195:100
  wire _col_2_n_u8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1194:100
  wire _col_2_d_x7_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1193:100
  wire _col_2_d_x7_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1193:100
  wire _col_2_d_x6_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1192:100
  wire _col_2_d_x6_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1192:100
  wire _col_2_d_x5_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1191:100
  wire _col_2_d_x5_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1191:100
  wire _col_2_d_x4_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1190:100
  wire _col_2_d_x4_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1190:100
  wire _col_2_d_x3_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1189:100
  wire _col_2_d_x3_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1189:100
  wire _col_2_d_x2_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1188:100
  wire _col_2_d_x2_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1188:100
  wire _col_2_d_x1_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1187:100
  wire _col_2_d_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1187:100
  wire _col_2_d_x0_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1186:100
  wire _col_2_d_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1186:100
  wire _col_2_n_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1185:100
  wire _col_2_n_t0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1184:83
  wire _col_2_n_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1183:83
  wire _col_2_n_w2_add_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1182:85
  wire _col_2_n_w2_sub_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1181:85
  wire _col_2_n_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1180:64
  wire _col_2_n_w3_add_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1179:85
  wire _col_2_n_w3_sub_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1178:85
  wire _col_2_n_w3_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1177:64
  wire _col_2_n_w1_add_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1176:85
  wire _col_2_n_w1_sub_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1175:85
  wire _col_2_n_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1174:64
  wire _col_2_n_c8192_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1173:73
  wire _col_2_n_c181_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1172:76
  wire _col_2_n_c181_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1171:76
  wire _col_2_n_c128_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1170:76
  wire _col_2_n_c128_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1169:76
  wire _col_2_n_c4_2_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1168:70
  wire _col_2_n_c4_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1167:70
  wire _col_2_n_c4_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1166:70
  wire _col_1_n_val_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1164:87
  wire _col_1_n_tmp_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1163:105
  wire _col_1_n_val_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1161:87
  wire _col_1_n_tmp_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1160:105
  wire _col_1_n_val_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1158:87
  wire _col_1_n_tmp_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1157:105
  wire _col_1_n_val_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1155:87
  wire _col_1_n_tmp_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1154:105
  wire _col_1_n_val_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1152:87
  wire _col_1_n_tmp_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1151:105
  wire _col_1_n_val_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1149:87
  wire _col_1_n_tmp_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1148:105
  wire _col_1_n_val_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1146:87
  wire _col_1_n_tmp_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1145:105
  wire _col_1_n_val_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1143:87
  wire _col_1_n_tmp_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1142:105
  wire _col_1_d_x4_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1141:100
  wire _col_1_d_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1141:100
  wire _col_1_n_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1140:83
  wire _col_1_n_w4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1139:100
  wire _col_1_n_v4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1138:100
  wire _col_1_n_u4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1137:100
  wire _col_1_d_x2_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1136:100
  wire _col_1_d_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1136:100
  wire _col_1_n_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1135:83
  wire _col_1_n_w2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1134:100
  wire _col_1_n_v2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1133:100
  wire _col_1_n_u2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1132:100
  wire _col_1_d_x0_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1131:100
  wire _col_1_d_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1131:100
  wire _col_1_n_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1130:100
  wire _col_1_d_x3_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1129:100
  wire _col_1_d_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1129:100
  wire _col_1_n_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1128:100
  wire _col_1_d_x8_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1127:100
  wire _col_1_d_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1127:100
  wire _col_1_n_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1126:100
  wire _col_1_d_x7_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1125:100
  wire _col_1_d_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1125:100
  wire _col_1_n_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1124:100
  wire _col_1_d_x5_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1123:100
  wire _col_1_d_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1123:100
  wire _col_1_n_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1122:100
  wire _col_1_d_x6_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1121:100
  wire _col_1_d_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1121:100
  wire _col_1_n_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1120:100
  wire _col_1_d_x4_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1119:100
  wire _col_1_d_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1119:100
  wire _col_1_n_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1118:100
  wire _col_1_d_x1_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1117:100
  wire _col_1_d_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1117:100
  wire _col_1_n_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1116:100
  wire _col_1_d_x3_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1115:100
  wire _col_1_d_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1115:100
  wire _col_1_n_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1114:83
  wire _col_1_n_v3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1113:100
  wire _col_1_n_u3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1112:100
  wire _col_1_d_x2_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1111:100
  wire _col_1_d_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1111:100
  wire _col_1_n_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1110:83
  wire _col_1_n_v2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1109:100
  wire _col_1_n_u2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1108:100
  wire _col_1_d_x1_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1107:100
  wire _col_1_d_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1107:100
  wire _col_1_n_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1106:100
  wire _col_1_n_v1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1105:100
  wire _col_1_n_u1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1104:100
  wire _col_1_d_x0_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1103:100
  wire _col_1_d_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1103:100
  wire _col_1_n_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1102:100
  wire _col_1_d_x8_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1101:100
  wire _col_1_d_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1101:100
  wire _col_1_n_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1100:100
  wire _col_1_d_x7_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1099:100
  wire _col_1_d_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1099:100
  wire _col_1_n_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1098:83
  wire _col_1_n_v7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1097:100
  wire _col_1_n_u7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1096:100
  wire _col_1_d_x6_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1095:100
  wire _col_1_d_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1095:100
  wire _col_1_n_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1094:83
  wire _col_1_n_v6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1093:100
  wire _col_1_n_u6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1092:100
  wire _col_1_d_x8_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1091:100
  wire _col_1_d_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1091:100
  wire _col_1_n_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1090:100
  wire _col_1_n_v8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1089:100
  wire _col_1_n_u8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1088:100
  wire _col_1_d_x5_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1087:100
  wire _col_1_d_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1087:100
  wire _col_1_n_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1086:83
  wire _col_1_n_v5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1085:100
  wire _col_1_n_u5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1084:100
  wire _col_1_d_x4_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1083:100
  wire _col_1_d_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1083:100
  wire _col_1_n_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1082:83
  wire _col_1_n_v4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1081:100
  wire _col_1_n_u4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1080:100
  wire _col_1_d_x8_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1079:100
  wire _col_1_d_x8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1079:100
  wire _col_1_n_x8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1078:100
  wire _col_1_n_v8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1077:100
  wire _col_1_n_u8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1076:100
  wire _col_1_d_x7_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1075:100
  wire _col_1_d_x7_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1075:100
  wire _col_1_d_x6_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1074:100
  wire _col_1_d_x6_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1074:100
  wire _col_1_d_x5_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1073:100
  wire _col_1_d_x5_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1073:100
  wire _col_1_d_x4_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1072:100
  wire _col_1_d_x4_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1072:100
  wire _col_1_d_x3_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1071:100
  wire _col_1_d_x3_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1071:100
  wire _col_1_d_x2_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1070:100
  wire _col_1_d_x2_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1070:100
  wire _col_1_d_x1_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1069:100
  wire _col_1_d_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1069:100
  wire _col_1_d_x0_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1068:100
  wire _col_1_d_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1068:100
  wire _col_1_n_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1067:100
  wire _col_1_n_t0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1066:83
  wire _col_1_n_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1065:83
  wire _col_1_n_w2_add_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1064:85
  wire _col_1_n_w2_sub_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1063:85
  wire _col_1_n_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1062:64
  wire _col_1_n_w3_add_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1061:85
  wire _col_1_n_w3_sub_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1060:85
  wire _col_1_n_w3_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1059:64
  wire _col_1_n_w1_add_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1058:85
  wire _col_1_n_w1_sub_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1057:85
  wire _col_1_n_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1056:64
  wire _col_1_n_c8192_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1055:73
  wire _col_1_n_c181_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1054:76
  wire _col_1_n_c181_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1053:76
  wire _col_1_n_c128_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1052:76
  wire _col_1_n_c128_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1051:76
  wire _col_1_n_c4_2_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1050:70
  wire _col_1_n_c4_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1049:70
  wire _col_1_n_c4_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1048:70
  wire _col_0_n_val_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1046:87
  wire _col_0_n_tmp_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1045:105
  wire _col_0_n_val_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1043:87
  wire _col_0_n_tmp_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1042:105
  wire _col_0_n_val_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1040:87
  wire _col_0_n_tmp_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1039:105
  wire _col_0_n_val_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1037:87
  wire _col_0_n_tmp_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1036:105
  wire _col_0_n_val_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1034:87
  wire _col_0_n_tmp_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1033:105
  wire _col_0_n_val_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1031:87
  wire _col_0_n_tmp_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1030:105
  wire _col_0_n_val_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1028:87
  wire _col_0_n_tmp_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1027:105
  wire _col_0_n_val_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1025:87
  wire _col_0_n_tmp_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1024:105
  wire _col_0_d_x4_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1023:100
  wire _col_0_d_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1023:100
  wire _col_0_n_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1022:83
  wire _col_0_n_w4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1021:100
  wire _col_0_n_v4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1020:100
  wire _col_0_n_u4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1019:100
  wire _col_0_d_x2_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1018:100
  wire _col_0_d_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1018:100
  wire _col_0_n_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1017:83
  wire _col_0_n_w2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1016:100
  wire _col_0_n_v2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1015:100
  wire _col_0_n_u2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1014:100
  wire _col_0_d_x0_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1013:100
  wire _col_0_d_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1013:100
  wire _col_0_n_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1012:100
  wire _col_0_d_x3_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1011:100
  wire _col_0_d_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1011:100
  wire _col_0_n_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1010:100
  wire _col_0_d_x8_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1009:100
  wire _col_0_d_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1009:100
  wire _col_0_n_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1008:100
  wire _col_0_d_x7_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1007:100
  wire _col_0_d_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1007:100
  wire _col_0_n_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1006:100
  wire _col_0_d_x5_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1005:100
  wire _col_0_d_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1005:100
  wire _col_0_n_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1004:100
  wire _col_0_d_x6_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1003:100
  wire _col_0_d_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1003:100
  wire _col_0_n_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1002:100
  wire _col_0_d_x4_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1001:100
  wire _col_0_d_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1001:100
  wire _col_0_n_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1000:100
  wire _col_0_d_x1_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:999:100
  wire _col_0_d_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:999:100
  wire _col_0_n_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:998:100
  wire _col_0_d_x3_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:997:100
  wire _col_0_d_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:997:100
  wire _col_0_n_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:996:83
  wire _col_0_n_v3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:995:100
  wire _col_0_n_u3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:994:100
  wire _col_0_d_x2_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:993:100
  wire _col_0_d_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:993:100
  wire _col_0_n_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:992:83
  wire _col_0_n_v2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:991:100
  wire _col_0_n_u2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:990:100
  wire _col_0_d_x1_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:989:100
  wire _col_0_d_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:989:100
  wire _col_0_n_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:988:100
  wire _col_0_n_v1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:987:100
  wire _col_0_n_u1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:986:100
  wire _col_0_d_x0_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:985:100
  wire _col_0_d_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:985:100
  wire _col_0_n_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:984:100
  wire _col_0_d_x8_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:983:100
  wire _col_0_d_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:983:100
  wire _col_0_n_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:982:100
  wire _col_0_d_x7_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:981:100
  wire _col_0_d_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:981:100
  wire _col_0_n_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:980:83
  wire _col_0_n_v7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:979:100
  wire _col_0_n_u7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:978:100
  wire _col_0_d_x6_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:977:100
  wire _col_0_d_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:977:100
  wire _col_0_n_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:976:83
  wire _col_0_n_v6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:975:100
  wire _col_0_n_u6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:974:100
  wire _col_0_d_x8_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:973:100
  wire _col_0_d_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:973:100
  wire _col_0_n_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:972:100
  wire _col_0_n_v8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:971:100
  wire _col_0_n_u8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:970:100
  wire _col_0_d_x5_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:969:100
  wire _col_0_d_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:969:100
  wire _col_0_n_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:968:83
  wire _col_0_n_v5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:967:100
  wire _col_0_n_u5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:966:100
  wire _col_0_d_x4_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:965:100
  wire _col_0_d_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:965:100
  wire _col_0_n_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:964:83
  wire _col_0_n_v4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:963:100
  wire _col_0_n_u4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:962:100
  wire _col_0_d_x8_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:961:100
  wire _col_0_d_x8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:961:100
  wire _col_0_n_x8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:960:100
  wire _col_0_n_v8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:959:100
  wire _col_0_n_u8_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:958:100
  wire _col_0_d_x7_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:957:100
  wire _col_0_d_x7_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:957:100
  wire _col_0_d_x6_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:956:100
  wire _col_0_d_x6_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:956:100
  wire _col_0_d_x5_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:955:100
  wire _col_0_d_x5_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:955:100
  wire _col_0_d_x4_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:954:100
  wire _col_0_d_x4_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:954:100
  wire _col_0_d_x3_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:953:100
  wire _col_0_d_x3_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:953:100
  wire _col_0_d_x2_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:952:100
  wire _col_0_d_x2_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:952:100
  wire _col_0_d_x1_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:951:100
  wire _col_0_d_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:951:100
  wire _col_0_d_x0_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:950:100
  wire _col_0_d_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:950:100
  wire _col_0_n_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:949:100
  wire _col_0_n_t0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:948:83
  wire _col_0_n_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:947:83
  wire _col_0_n_w2_add_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:946:85
  wire _col_0_n_w2_sub_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:945:85
  wire _col_0_n_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:944:64
  wire _col_0_n_w3_add_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:943:85
  wire _col_0_n_w3_sub_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:942:85
  wire _col_0_n_w3_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:941:64
  wire _col_0_n_w1_add_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:940:85
  wire _col_0_n_w1_sub_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:939:85
  wire _col_0_n_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:938:64
  wire _col_0_n_c8192_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:937:73
  wire _col_0_n_c181_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:936:76
  wire _col_0_n_c181_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:935:76
  wire _col_0_n_c128_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:934:76
  wire _col_0_n_c128_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:933:76
  wire _col_0_n_c4_2_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:932:70
  wire _col_0_n_c4_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:931:70
  wire _col_0_n_c4_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:930:70
  wire _row_7_n_shr_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:929:87
  wire _row_7_n_tmp_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:928:105
  wire _row_7_n_shr_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:927:87
  wire _row_7_n_tmp_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:926:105
  wire _row_7_n_shr_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:925:87
  wire _row_7_n_tmp_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:924:105
  wire _row_7_n_shr_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:923:87
  wire _row_7_n_tmp_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:922:105
  wire _row_7_n_shr_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:921:87
  wire _row_7_n_tmp_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:920:105
  wire _row_7_n_shr_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:919:87
  wire _row_7_n_tmp_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:918:105
  wire _row_7_n_shr_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:917:87
  wire _row_7_n_tmp_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:916:105
  wire _row_7_n_shr_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:915:87
  wire _row_7_n_tmp_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:914:105
  wire _row_7_d_x4_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:913:100
  wire _row_7_d_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:913:100
  wire _row_7_n_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:912:83
  wire _row_7_n_w4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:911:100
  wire _row_7_n_v4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:910:100
  wire _row_7_n_u4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:909:100
  wire _row_7_d_x2_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:908:100
  wire _row_7_d_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:908:100
  wire _row_7_n_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:907:83
  wire _row_7_n_w2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:906:100
  wire _row_7_n_v2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:905:100
  wire _row_7_n_u2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:904:100
  wire _row_7_d_x0_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:903:100
  wire _row_7_d_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:903:100
  wire _row_7_n_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:902:100
  wire _row_7_d_x3_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:901:100
  wire _row_7_d_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:901:100
  wire _row_7_n_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:900:100
  wire _row_7_d_x8_4_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:899:100
  wire _row_7_d_x8_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:899:100
  wire _row_7_n_x8_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:898:100
  wire _row_7_d_x7_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:897:100
  wire _row_7_d_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:897:100
  wire _row_7_n_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:896:100
  wire _row_7_d_x5_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:895:100
  wire _row_7_d_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:895:100
  wire _row_7_n_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:894:100
  wire _row_7_d_x6_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:893:100
  wire _row_7_d_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:893:100
  wire _row_7_n_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:892:100
  wire _row_7_d_x4_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:891:100
  wire _row_7_d_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:891:100
  wire _row_7_n_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:890:100
  wire _row_7_d_x1_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:889:100
  wire _row_7_d_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:889:100
  wire _row_7_n_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:888:100
  wire _row_7_d_x3_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:887:100
  wire _row_7_d_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:887:100
  wire _row_7_n_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:886:100
  wire _row_7_n_t3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:885:100
  wire _row_7_d_x2_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:884:100
  wire _row_7_d_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:884:100
  wire _row_7_n_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:883:100
  wire _row_7_n_t2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:882:100
  wire _row_7_d_x1_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:881:100
  wire _row_7_d_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:881:100
  wire _row_7_n_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:880:100
  wire _row_7_n_t1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:879:100
  wire _row_7_d_x0_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:878:100
  wire _row_7_d_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:878:100
  wire _row_7_n_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:877:100
  wire _row_7_d_x8_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:876:100
  wire _row_7_d_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:876:100
  wire _row_7_n_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:875:100
  wire _row_7_d_x7_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:874:100
  wire _row_7_d_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:874:100
  wire _row_7_n_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:873:100
  wire _row_7_n_t7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:872:100
  wire _row_7_d_x6_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:871:100
  wire _row_7_d_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:871:100
  wire _row_7_n_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:870:100
  wire _row_7_n_t6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:869:100
  wire _row_7_d_x8_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:868:100
  wire _row_7_d_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:868:100
  wire _row_7_n_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:867:100
  wire _row_7_n_t8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:866:100
  wire _row_7_d_x5_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:865:100
  wire _row_7_d_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:865:100
  wire _row_7_n_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:864:100
  wire _row_7_n_t5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:863:100
  wire _row_7_d_x4_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:862:100
  wire _row_7_d_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:862:100
  wire _row_7_n_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:861:100
  wire _row_7_n_t4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:860:100
  wire _row_7_d_x8_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:859:100
  wire _row_7_d_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:859:100
  wire _row_7_n_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:858:100
  wire _row_7_n_t8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:857:100
  wire _row_7_d_x7_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:856:100
  wire _row_7_d_x7_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:856:100
  wire _row_7_d_x6_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:855:100
  wire _row_7_d_x6_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:855:100
  wire _row_7_d_x5_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:854:100
  wire _row_7_d_x5_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:854:100
  wire _row_7_d_x4_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:853:100
  wire _row_7_d_x4_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:853:100
  wire _row_7_d_x3_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:852:100
  wire _row_7_d_x3_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:852:100
  wire _row_7_d_x2_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:851:100
  wire _row_7_d_x2_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:851:100
  wire _row_7_d_x1_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:850:100
  wire _row_7_d_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:850:100
  wire _row_7_d_x0_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:849:100
  wire _row_7_d_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:849:100
  wire _row_7_n_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:848:100
  wire _row_7_n_t0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:847:83
  wire _row_7_n_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:846:83
  wire _row_7_n_w2_add_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:845:85
  wire _row_7_n_w2_sub_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:844:85
  wire _row_7_n_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:843:64
  wire _row_7_n_w3_add_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:842:85
  wire _row_7_n_w3_sub_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:841:85
  wire _row_7_n_w3_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:840:64
  wire _row_7_n_w1_add_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:839:85
  wire _row_7_n_w1_sub_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:838:85
  wire _row_7_n_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:837:64
  wire _row_7_n_c181_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:836:76
  wire _row_7_n_c181_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:835:76
  wire _row_7_n_c128_2_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:834:76
  wire _row_7_n_c128_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:833:76
  wire _row_7_n_c128_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:832:76
  wire _row_6_n_shr_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:831:87
  wire _row_6_n_tmp_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:830:105
  wire _row_6_n_shr_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:829:87
  wire _row_6_n_tmp_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:828:105
  wire _row_6_n_shr_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:827:87
  wire _row_6_n_tmp_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:826:105
  wire _row_6_n_shr_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:825:87
  wire _row_6_n_tmp_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:824:105
  wire _row_6_n_shr_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:823:87
  wire _row_6_n_tmp_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:822:105
  wire _row_6_n_shr_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:821:87
  wire _row_6_n_tmp_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:820:105
  wire _row_6_n_shr_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:819:87
  wire _row_6_n_tmp_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:818:105
  wire _row_6_n_shr_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:817:87
  wire _row_6_n_tmp_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:816:105
  wire _row_6_d_x4_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:815:100
  wire _row_6_d_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:815:100
  wire _row_6_n_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:814:83
  wire _row_6_n_w4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:813:100
  wire _row_6_n_v4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:812:100
  wire _row_6_n_u4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:811:100
  wire _row_6_d_x2_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:810:100
  wire _row_6_d_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:810:100
  wire _row_6_n_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:809:83
  wire _row_6_n_w2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:808:100
  wire _row_6_n_v2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:807:100
  wire _row_6_n_u2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:806:100
  wire _row_6_d_x0_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:805:100
  wire _row_6_d_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:805:100
  wire _row_6_n_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:804:100
  wire _row_6_d_x3_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:803:100
  wire _row_6_d_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:803:100
  wire _row_6_n_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:802:100
  wire _row_6_d_x8_4_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:801:100
  wire _row_6_d_x8_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:801:100
  wire _row_6_n_x8_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:800:100
  wire _row_6_d_x7_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:799:100
  wire _row_6_d_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:799:100
  wire _row_6_n_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:798:100
  wire _row_6_d_x5_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:797:100
  wire _row_6_d_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:797:100
  wire _row_6_n_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:796:100
  wire _row_6_d_x6_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:795:100
  wire _row_6_d_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:795:100
  wire _row_6_n_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:794:100
  wire _row_6_d_x4_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:793:100
  wire _row_6_d_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:793:100
  wire _row_6_n_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:792:100
  wire _row_6_d_x1_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:791:100
  wire _row_6_d_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:791:100
  wire _row_6_n_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:790:100
  wire _row_6_d_x3_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:789:100
  wire _row_6_d_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:789:100
  wire _row_6_n_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:788:100
  wire _row_6_n_t3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:787:100
  wire _row_6_d_x2_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:786:100
  wire _row_6_d_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:786:100
  wire _row_6_n_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:785:100
  wire _row_6_n_t2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:784:100
  wire _row_6_d_x1_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:783:100
  wire _row_6_d_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:783:100
  wire _row_6_n_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:782:100
  wire _row_6_n_t1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:781:100
  wire _row_6_d_x0_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:780:100
  wire _row_6_d_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:780:100
  wire _row_6_n_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:779:100
  wire _row_6_d_x8_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:778:100
  wire _row_6_d_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:778:100
  wire _row_6_n_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:777:100
  wire _row_6_d_x7_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:776:100
  wire _row_6_d_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:776:100
  wire _row_6_n_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:775:100
  wire _row_6_n_t7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:774:100
  wire _row_6_d_x6_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:773:100
  wire _row_6_d_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:773:100
  wire _row_6_n_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:772:100
  wire _row_6_n_t6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:771:100
  wire _row_6_d_x8_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:770:100
  wire _row_6_d_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:770:100
  wire _row_6_n_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:769:100
  wire _row_6_n_t8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:768:100
  wire _row_6_d_x5_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:767:100
  wire _row_6_d_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:767:100
  wire _row_6_n_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:766:100
  wire _row_6_n_t5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:765:100
  wire _row_6_d_x4_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:764:100
  wire _row_6_d_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:764:100
  wire _row_6_n_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:763:100
  wire _row_6_n_t4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:762:100
  wire _row_6_d_x8_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:761:100
  wire _row_6_d_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:761:100
  wire _row_6_n_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:760:100
  wire _row_6_n_t8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:759:100
  wire _row_6_d_x7_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:758:100
  wire _row_6_d_x7_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:758:100
  wire _row_6_d_x6_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:757:100
  wire _row_6_d_x6_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:757:100
  wire _row_6_d_x5_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:756:100
  wire _row_6_d_x5_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:756:100
  wire _row_6_d_x4_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:755:100
  wire _row_6_d_x4_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:755:100
  wire _row_6_d_x3_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:754:100
  wire _row_6_d_x3_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:754:100
  wire _row_6_d_x2_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:753:100
  wire _row_6_d_x2_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:753:100
  wire _row_6_d_x1_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:752:100
  wire _row_6_d_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:752:100
  wire _row_6_d_x0_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:751:100
  wire _row_6_d_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:751:100
  wire _row_6_n_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:750:100
  wire _row_6_n_t0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:749:83
  wire _row_6_n_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:748:83
  wire _row_6_n_w2_add_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:747:85
  wire _row_6_n_w2_sub_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:746:85
  wire _row_6_n_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:745:64
  wire _row_6_n_w3_add_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:744:85
  wire _row_6_n_w3_sub_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:743:85
  wire _row_6_n_w3_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:742:64
  wire _row_6_n_w1_add_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:741:85
  wire _row_6_n_w1_sub_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:740:85
  wire _row_6_n_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:739:64
  wire _row_6_n_c181_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:738:76
  wire _row_6_n_c181_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:737:76
  wire _row_6_n_c128_2_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:736:76
  wire _row_6_n_c128_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:735:76
  wire _row_6_n_c128_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:734:76
  wire _row_5_n_shr_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:733:87
  wire _row_5_n_tmp_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:732:105
  wire _row_5_n_shr_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:731:87
  wire _row_5_n_tmp_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:730:105
  wire _row_5_n_shr_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:729:87
  wire _row_5_n_tmp_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:728:105
  wire _row_5_n_shr_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:727:87
  wire _row_5_n_tmp_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:726:105
  wire _row_5_n_shr_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:725:87
  wire _row_5_n_tmp_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:724:105
  wire _row_5_n_shr_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:723:87
  wire _row_5_n_tmp_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:722:105
  wire _row_5_n_shr_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:721:87
  wire _row_5_n_tmp_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:720:105
  wire _row_5_n_shr_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:719:87
  wire _row_5_n_tmp_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:718:105
  wire _row_5_d_x4_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:717:100
  wire _row_5_d_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:717:100
  wire _row_5_n_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:716:83
  wire _row_5_n_w4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:715:100
  wire _row_5_n_v4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:714:100
  wire _row_5_n_u4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:713:100
  wire _row_5_d_x2_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:712:100
  wire _row_5_d_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:712:100
  wire _row_5_n_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:711:83
  wire _row_5_n_w2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:710:100
  wire _row_5_n_v2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:709:100
  wire _row_5_n_u2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:708:100
  wire _row_5_d_x0_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:707:100
  wire _row_5_d_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:707:100
  wire _row_5_n_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:706:100
  wire _row_5_d_x3_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:705:100
  wire _row_5_d_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:705:100
  wire _row_5_n_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:704:100
  wire _row_5_d_x8_4_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:703:100
  wire _row_5_d_x8_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:703:100
  wire _row_5_n_x8_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:702:100
  wire _row_5_d_x7_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:701:100
  wire _row_5_d_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:701:100
  wire _row_5_n_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:700:100
  wire _row_5_d_x5_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:699:100
  wire _row_5_d_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:699:100
  wire _row_5_n_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:698:100
  wire _row_5_d_x6_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:697:100
  wire _row_5_d_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:697:100
  wire _row_5_n_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:696:100
  wire _row_5_d_x4_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:695:100
  wire _row_5_d_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:695:100
  wire _row_5_n_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:694:100
  wire _row_5_d_x1_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:693:100
  wire _row_5_d_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:693:100
  wire _row_5_n_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:692:100
  wire _row_5_d_x3_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:691:100
  wire _row_5_d_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:691:100
  wire _row_5_n_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:690:100
  wire _row_5_n_t3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:689:100
  wire _row_5_d_x2_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:688:100
  wire _row_5_d_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:688:100
  wire _row_5_n_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:687:100
  wire _row_5_n_t2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:686:100
  wire _row_5_d_x1_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:685:100
  wire _row_5_d_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:685:100
  wire _row_5_n_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:684:100
  wire _row_5_n_t1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:683:100
  wire _row_5_d_x0_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:682:100
  wire _row_5_d_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:682:100
  wire _row_5_n_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:681:100
  wire _row_5_d_x8_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:680:100
  wire _row_5_d_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:680:100
  wire _row_5_n_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:679:100
  wire _row_5_d_x7_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:678:100
  wire _row_5_d_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:678:100
  wire _row_5_n_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:677:100
  wire _row_5_n_t7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:676:100
  wire _row_5_d_x6_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:675:100
  wire _row_5_d_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:675:100
  wire _row_5_n_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:674:100
  wire _row_5_n_t6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:673:100
  wire _row_5_d_x8_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:672:100
  wire _row_5_d_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:672:100
  wire _row_5_n_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:671:100
  wire _row_5_n_t8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:670:100
  wire _row_5_d_x5_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:669:100
  wire _row_5_d_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:669:100
  wire _row_5_n_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:668:100
  wire _row_5_n_t5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:667:100
  wire _row_5_d_x4_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:666:100
  wire _row_5_d_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:666:100
  wire _row_5_n_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:665:100
  wire _row_5_n_t4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:664:100
  wire _row_5_d_x8_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:663:100
  wire _row_5_d_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:663:100
  wire _row_5_n_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:662:100
  wire _row_5_n_t8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:661:100
  wire _row_5_d_x7_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:660:100
  wire _row_5_d_x7_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:660:100
  wire _row_5_d_x6_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:659:100
  wire _row_5_d_x6_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:659:100
  wire _row_5_d_x5_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:658:100
  wire _row_5_d_x5_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:658:100
  wire _row_5_d_x4_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:657:100
  wire _row_5_d_x4_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:657:100
  wire _row_5_d_x3_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:656:100
  wire _row_5_d_x3_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:656:100
  wire _row_5_d_x2_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:655:100
  wire _row_5_d_x2_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:655:100
  wire _row_5_d_x1_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:654:100
  wire _row_5_d_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:654:100
  wire _row_5_d_x0_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:653:100
  wire _row_5_d_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:653:100
  wire _row_5_n_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:652:100
  wire _row_5_n_t0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:651:83
  wire _row_5_n_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:650:83
  wire _row_5_n_w2_add_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:649:85
  wire _row_5_n_w2_sub_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:648:85
  wire _row_5_n_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:647:64
  wire _row_5_n_w3_add_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:646:85
  wire _row_5_n_w3_sub_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:645:85
  wire _row_5_n_w3_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:644:64
  wire _row_5_n_w1_add_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:643:85
  wire _row_5_n_w1_sub_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:642:85
  wire _row_5_n_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:641:64
  wire _row_5_n_c181_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:640:76
  wire _row_5_n_c181_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:639:76
  wire _row_5_n_c128_2_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:638:76
  wire _row_5_n_c128_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:637:76
  wire _row_5_n_c128_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:636:76
  wire _row_4_n_shr_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:635:87
  wire _row_4_n_tmp_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:634:105
  wire _row_4_n_shr_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:633:87
  wire _row_4_n_tmp_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:632:105
  wire _row_4_n_shr_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:631:87
  wire _row_4_n_tmp_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:630:105
  wire _row_4_n_shr_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:629:87
  wire _row_4_n_tmp_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:628:105
  wire _row_4_n_shr_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:627:87
  wire _row_4_n_tmp_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:626:105
  wire _row_4_n_shr_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:625:87
  wire _row_4_n_tmp_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:624:105
  wire _row_4_n_shr_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:623:87
  wire _row_4_n_tmp_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:622:105
  wire _row_4_n_shr_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:621:87
  wire _row_4_n_tmp_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:620:105
  wire _row_4_d_x4_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:619:100
  wire _row_4_d_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:619:100
  wire _row_4_n_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:618:83
  wire _row_4_n_w4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:617:100
  wire _row_4_n_v4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:616:100
  wire _row_4_n_u4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:615:100
  wire _row_4_d_x2_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:614:100
  wire _row_4_d_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:614:100
  wire _row_4_n_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:613:83
  wire _row_4_n_w2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:612:100
  wire _row_4_n_v2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:611:100
  wire _row_4_n_u2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:610:100
  wire _row_4_d_x0_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:609:100
  wire _row_4_d_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:609:100
  wire _row_4_n_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:608:100
  wire _row_4_d_x3_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:607:100
  wire _row_4_d_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:607:100
  wire _row_4_n_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:606:100
  wire _row_4_d_x8_4_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:605:100
  wire _row_4_d_x8_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:605:100
  wire _row_4_n_x8_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:604:100
  wire _row_4_d_x7_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:603:100
  wire _row_4_d_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:603:100
  wire _row_4_n_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:602:100
  wire _row_4_d_x5_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:601:100
  wire _row_4_d_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:601:100
  wire _row_4_n_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:600:100
  wire _row_4_d_x6_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:599:100
  wire _row_4_d_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:599:100
  wire _row_4_n_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:598:100
  wire _row_4_d_x4_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:597:100
  wire _row_4_d_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:597:100
  wire _row_4_n_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:596:100
  wire _row_4_d_x1_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:595:100
  wire _row_4_d_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:595:100
  wire _row_4_n_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:594:100
  wire _row_4_d_x3_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:593:100
  wire _row_4_d_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:593:100
  wire _row_4_n_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:592:100
  wire _row_4_n_t3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:591:100
  wire _row_4_d_x2_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:590:100
  wire _row_4_d_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:590:100
  wire _row_4_n_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:589:100
  wire _row_4_n_t2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:588:100
  wire _row_4_d_x1_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:587:100
  wire _row_4_d_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:587:100
  wire _row_4_n_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:586:100
  wire _row_4_n_t1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:585:100
  wire _row_4_d_x0_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:584:100
  wire _row_4_d_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:584:100
  wire _row_4_n_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:583:100
  wire _row_4_d_x8_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:582:100
  wire _row_4_d_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:582:100
  wire _row_4_n_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:581:100
  wire _row_4_d_x7_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:580:100
  wire _row_4_d_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:580:100
  wire _row_4_n_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:579:100
  wire _row_4_n_t7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:578:100
  wire _row_4_d_x6_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:577:100
  wire _row_4_d_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:577:100
  wire _row_4_n_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:576:100
  wire _row_4_n_t6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:575:100
  wire _row_4_d_x8_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:574:100
  wire _row_4_d_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:574:100
  wire _row_4_n_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:573:100
  wire _row_4_n_t8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:572:100
  wire _row_4_d_x5_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:571:100
  wire _row_4_d_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:571:100
  wire _row_4_n_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:570:100
  wire _row_4_n_t5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:569:100
  wire _row_4_d_x4_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:568:100
  wire _row_4_d_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:568:100
  wire _row_4_n_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:567:100
  wire _row_4_n_t4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:566:100
  wire _row_4_d_x8_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:565:100
  wire _row_4_d_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:565:100
  wire _row_4_n_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:564:100
  wire _row_4_n_t8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:563:100
  wire _row_4_d_x7_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:562:100
  wire _row_4_d_x7_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:562:100
  wire _row_4_d_x6_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:561:100
  wire _row_4_d_x6_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:561:100
  wire _row_4_d_x5_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:560:100
  wire _row_4_d_x5_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:560:100
  wire _row_4_d_x4_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:559:100
  wire _row_4_d_x4_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:559:100
  wire _row_4_d_x3_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:558:100
  wire _row_4_d_x3_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:558:100
  wire _row_4_d_x2_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:557:100
  wire _row_4_d_x2_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:557:100
  wire _row_4_d_x1_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:556:100
  wire _row_4_d_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:556:100
  wire _row_4_d_x0_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:555:100
  wire _row_4_d_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:555:100
  wire _row_4_n_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:554:100
  wire _row_4_n_t0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:553:83
  wire _row_4_n_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:552:83
  wire _row_4_n_w2_add_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:551:85
  wire _row_4_n_w2_sub_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:550:85
  wire _row_4_n_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:549:64
  wire _row_4_n_w3_add_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:548:85
  wire _row_4_n_w3_sub_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:547:85
  wire _row_4_n_w3_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:546:64
  wire _row_4_n_w1_add_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:545:85
  wire _row_4_n_w1_sub_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:544:85
  wire _row_4_n_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:543:64
  wire _row_4_n_c181_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:542:76
  wire _row_4_n_c181_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:541:76
  wire _row_4_n_c128_2_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:540:76
  wire _row_4_n_c128_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:539:76
  wire _row_4_n_c128_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:538:76
  wire _row_3_n_shr_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:537:87
  wire _row_3_n_tmp_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:536:105
  wire _row_3_n_shr_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:535:87
  wire _row_3_n_tmp_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:534:105
  wire _row_3_n_shr_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:533:87
  wire _row_3_n_tmp_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:532:105
  wire _row_3_n_shr_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:531:87
  wire _row_3_n_tmp_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:530:105
  wire _row_3_n_shr_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:529:87
  wire _row_3_n_tmp_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:528:105
  wire _row_3_n_shr_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:527:87
  wire _row_3_n_tmp_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:526:105
  wire _row_3_n_shr_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:525:87
  wire _row_3_n_tmp_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:524:105
  wire _row_3_n_shr_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:523:87
  wire _row_3_n_tmp_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:522:105
  wire _row_3_d_x4_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:521:100
  wire _row_3_d_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:521:100
  wire _row_3_n_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:520:83
  wire _row_3_n_w4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:519:100
  wire _row_3_n_v4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:518:100
  wire _row_3_n_u4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:517:100
  wire _row_3_d_x2_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:516:100
  wire _row_3_d_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:516:100
  wire _row_3_n_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:515:83
  wire _row_3_n_w2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:514:100
  wire _row_3_n_v2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:513:100
  wire _row_3_n_u2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:512:100
  wire _row_3_d_x0_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:511:100
  wire _row_3_d_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:511:100
  wire _row_3_n_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:510:100
  wire _row_3_d_x3_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:509:100
  wire _row_3_d_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:509:100
  wire _row_3_n_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:508:100
  wire _row_3_d_x8_4_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:507:100
  wire _row_3_d_x8_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:507:100
  wire _row_3_n_x8_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:506:100
  wire _row_3_d_x7_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:505:100
  wire _row_3_d_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:505:100
  wire _row_3_n_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:504:100
  wire _row_3_d_x5_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:503:100
  wire _row_3_d_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:503:100
  wire _row_3_n_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:502:100
  wire _row_3_d_x6_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:501:100
  wire _row_3_d_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:501:100
  wire _row_3_n_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:500:100
  wire _row_3_d_x4_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:499:100
  wire _row_3_d_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:499:100
  wire _row_3_n_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:498:100
  wire _row_3_d_x1_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:497:100
  wire _row_3_d_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:497:100
  wire _row_3_n_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:496:100
  wire _row_3_d_x3_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:495:100
  wire _row_3_d_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:495:100
  wire _row_3_n_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:494:100
  wire _row_3_n_t3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:493:100
  wire _row_3_d_x2_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:492:100
  wire _row_3_d_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:492:100
  wire _row_3_n_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:491:100
  wire _row_3_n_t2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:490:100
  wire _row_3_d_x1_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:489:100
  wire _row_3_d_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:489:100
  wire _row_3_n_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:488:100
  wire _row_3_n_t1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:487:100
  wire _row_3_d_x0_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:486:100
  wire _row_3_d_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:486:100
  wire _row_3_n_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:485:100
  wire _row_3_d_x8_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:484:100
  wire _row_3_d_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:484:100
  wire _row_3_n_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:483:100
  wire _row_3_d_x7_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:482:100
  wire _row_3_d_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:482:100
  wire _row_3_n_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:481:100
  wire _row_3_n_t7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:480:100
  wire _row_3_d_x6_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:479:100
  wire _row_3_d_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:479:100
  wire _row_3_n_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:478:100
  wire _row_3_n_t6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:477:100
  wire _row_3_d_x8_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:476:100
  wire _row_3_d_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:476:100
  wire _row_3_n_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:475:100
  wire _row_3_n_t8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:474:100
  wire _row_3_d_x5_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:473:100
  wire _row_3_d_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:473:100
  wire _row_3_n_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:472:100
  wire _row_3_n_t5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:471:100
  wire _row_3_d_x4_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:470:100
  wire _row_3_d_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:470:100
  wire _row_3_n_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:469:100
  wire _row_3_n_t4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:468:100
  wire _row_3_d_x8_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:467:100
  wire _row_3_d_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:467:100
  wire _row_3_n_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:466:100
  wire _row_3_n_t8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:465:100
  wire _row_3_d_x7_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:464:100
  wire _row_3_d_x7_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:464:100
  wire _row_3_d_x6_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:463:100
  wire _row_3_d_x6_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:463:100
  wire _row_3_d_x5_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:462:100
  wire _row_3_d_x5_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:462:100
  wire _row_3_d_x4_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:461:100
  wire _row_3_d_x4_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:461:100
  wire _row_3_d_x3_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:460:100
  wire _row_3_d_x3_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:460:100
  wire _row_3_d_x2_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:459:100
  wire _row_3_d_x2_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:459:100
  wire _row_3_d_x1_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:458:100
  wire _row_3_d_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:458:100
  wire _row_3_d_x0_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:457:100
  wire _row_3_d_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:457:100
  wire _row_3_n_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:456:100
  wire _row_3_n_t0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:455:83
  wire _row_3_n_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:454:83
  wire _row_3_n_w2_add_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:453:85
  wire _row_3_n_w2_sub_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:452:85
  wire _row_3_n_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:451:64
  wire _row_3_n_w3_add_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:450:85
  wire _row_3_n_w3_sub_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:449:85
  wire _row_3_n_w3_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:448:64
  wire _row_3_n_w1_add_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:447:85
  wire _row_3_n_w1_sub_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:446:85
  wire _row_3_n_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:445:64
  wire _row_3_n_c181_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:444:76
  wire _row_3_n_c181_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:443:76
  wire _row_3_n_c128_2_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:442:76
  wire _row_3_n_c128_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:441:76
  wire _row_3_n_c128_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:440:76
  wire _row_2_n_shr_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:439:87
  wire _row_2_n_tmp_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:438:105
  wire _row_2_n_shr_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:437:87
  wire _row_2_n_tmp_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:436:105
  wire _row_2_n_shr_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:435:87
  wire _row_2_n_tmp_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:434:105
  wire _row_2_n_shr_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:433:87
  wire _row_2_n_tmp_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:432:105
  wire _row_2_n_shr_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:431:87
  wire _row_2_n_tmp_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:430:105
  wire _row_2_n_shr_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:429:87
  wire _row_2_n_tmp_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:428:105
  wire _row_2_n_shr_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:427:87
  wire _row_2_n_tmp_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:426:105
  wire _row_2_n_shr_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:425:87
  wire _row_2_n_tmp_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:424:105
  wire _row_2_d_x4_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:423:100
  wire _row_2_d_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:423:100
  wire _row_2_n_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:422:83
  wire _row_2_n_w4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:421:100
  wire _row_2_n_v4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:420:100
  wire _row_2_n_u4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:419:100
  wire _row_2_d_x2_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:418:100
  wire _row_2_d_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:418:100
  wire _row_2_n_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:417:83
  wire _row_2_n_w2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:416:100
  wire _row_2_n_v2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:415:100
  wire _row_2_n_u2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:414:100
  wire _row_2_d_x0_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:413:100
  wire _row_2_d_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:413:100
  wire _row_2_n_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:412:100
  wire _row_2_d_x3_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:411:100
  wire _row_2_d_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:411:100
  wire _row_2_n_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:410:100
  wire _row_2_d_x8_4_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:409:100
  wire _row_2_d_x8_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:409:100
  wire _row_2_n_x8_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:408:100
  wire _row_2_d_x7_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:407:100
  wire _row_2_d_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:407:100
  wire _row_2_n_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:406:100
  wire _row_2_d_x5_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:405:100
  wire _row_2_d_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:405:100
  wire _row_2_n_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:404:100
  wire _row_2_d_x6_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:403:100
  wire _row_2_d_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:403:100
  wire _row_2_n_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:402:100
  wire _row_2_d_x4_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:401:100
  wire _row_2_d_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:401:100
  wire _row_2_n_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:400:100
  wire _row_2_d_x1_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:399:100
  wire _row_2_d_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:399:100
  wire _row_2_n_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:398:100
  wire _row_2_d_x3_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:397:100
  wire _row_2_d_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:397:100
  wire _row_2_n_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:396:100
  wire _row_2_n_t3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:395:100
  wire _row_2_d_x2_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:394:100
  wire _row_2_d_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:394:100
  wire _row_2_n_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:393:100
  wire _row_2_n_t2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:392:100
  wire _row_2_d_x1_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:391:100
  wire _row_2_d_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:391:100
  wire _row_2_n_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:390:100
  wire _row_2_n_t1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:389:100
  wire _row_2_d_x0_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:388:100
  wire _row_2_d_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:388:100
  wire _row_2_n_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:387:100
  wire _row_2_d_x8_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:386:100
  wire _row_2_d_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:386:100
  wire _row_2_n_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:385:100
  wire _row_2_d_x7_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:384:100
  wire _row_2_d_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:384:100
  wire _row_2_n_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:383:100
  wire _row_2_n_t7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:382:100
  wire _row_2_d_x6_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:381:100
  wire _row_2_d_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:381:100
  wire _row_2_n_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:380:100
  wire _row_2_n_t6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:379:100
  wire _row_2_d_x8_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:378:100
  wire _row_2_d_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:378:100
  wire _row_2_n_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:377:100
  wire _row_2_n_t8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:376:100
  wire _row_2_d_x5_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:375:100
  wire _row_2_d_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:375:100
  wire _row_2_n_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:374:100
  wire _row_2_n_t5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:373:100
  wire _row_2_d_x4_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:372:100
  wire _row_2_d_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:372:100
  wire _row_2_n_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:371:100
  wire _row_2_n_t4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:370:100
  wire _row_2_d_x8_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:369:100
  wire _row_2_d_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:369:100
  wire _row_2_n_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:368:100
  wire _row_2_n_t8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:367:100
  wire _row_2_d_x7_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:366:100
  wire _row_2_d_x7_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:366:100
  wire _row_2_d_x6_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:365:100
  wire _row_2_d_x6_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:365:100
  wire _row_2_d_x5_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:364:100
  wire _row_2_d_x5_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:364:100
  wire _row_2_d_x4_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:363:100
  wire _row_2_d_x4_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:363:100
  wire _row_2_d_x3_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:362:100
  wire _row_2_d_x3_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:362:100
  wire _row_2_d_x2_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:361:100
  wire _row_2_d_x2_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:361:100
  wire _row_2_d_x1_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:360:100
  wire _row_2_d_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:360:100
  wire _row_2_d_x0_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:359:100
  wire _row_2_d_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:359:100
  wire _row_2_n_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:358:100
  wire _row_2_n_t0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:357:83
  wire _row_2_n_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:356:83
  wire _row_2_n_w2_add_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:355:85
  wire _row_2_n_w2_sub_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:354:85
  wire _row_2_n_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:353:64
  wire _row_2_n_w3_add_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:352:85
  wire _row_2_n_w3_sub_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:351:85
  wire _row_2_n_w3_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:350:64
  wire _row_2_n_w1_add_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:349:85
  wire _row_2_n_w1_sub_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:348:85
  wire _row_2_n_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:347:64
  wire _row_2_n_c181_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:346:76
  wire _row_2_n_c181_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:345:76
  wire _row_2_n_c128_2_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:344:76
  wire _row_2_n_c128_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:343:76
  wire _row_2_n_c128_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:342:76
  wire _row_1_n_shr_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:341:87
  wire _row_1_n_tmp_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:340:105
  wire _row_1_n_shr_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:339:87
  wire _row_1_n_tmp_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:338:105
  wire _row_1_n_shr_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:337:87
  wire _row_1_n_tmp_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:336:105
  wire _row_1_n_shr_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:335:87
  wire _row_1_n_tmp_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:334:105
  wire _row_1_n_shr_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:333:87
  wire _row_1_n_tmp_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:332:105
  wire _row_1_n_shr_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:331:87
  wire _row_1_n_tmp_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:330:105
  wire _row_1_n_shr_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:329:87
  wire _row_1_n_tmp_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:328:105
  wire _row_1_n_shr_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:327:87
  wire _row_1_n_tmp_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:326:105
  wire _row_1_d_x4_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:325:100
  wire _row_1_d_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:325:100
  wire _row_1_n_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:324:83
  wire _row_1_n_w4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:323:100
  wire _row_1_n_v4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:322:100
  wire _row_1_n_u4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:321:100
  wire _row_1_d_x2_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:320:100
  wire _row_1_d_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:320:100
  wire _row_1_n_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:319:83
  wire _row_1_n_w2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:318:100
  wire _row_1_n_v2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:317:100
  wire _row_1_n_u2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:316:100
  wire _row_1_d_x0_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:315:100
  wire _row_1_d_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:315:100
  wire _row_1_n_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:314:100
  wire _row_1_d_x3_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:313:100
  wire _row_1_d_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:313:100
  wire _row_1_n_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:312:100
  wire _row_1_d_x8_4_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:311:100
  wire _row_1_d_x8_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:311:100
  wire _row_1_n_x8_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:310:100
  wire _row_1_d_x7_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:309:100
  wire _row_1_d_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:309:100
  wire _row_1_n_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:308:100
  wire _row_1_d_x5_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:307:100
  wire _row_1_d_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:307:100
  wire _row_1_n_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:306:100
  wire _row_1_d_x6_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:305:100
  wire _row_1_d_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:305:100
  wire _row_1_n_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:304:100
  wire _row_1_d_x4_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:303:100
  wire _row_1_d_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:303:100
  wire _row_1_n_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:302:100
  wire _row_1_d_x1_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:301:100
  wire _row_1_d_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:301:100
  wire _row_1_n_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:300:100
  wire _row_1_d_x3_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:299:100
  wire _row_1_d_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:299:100
  wire _row_1_n_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:298:100
  wire _row_1_n_t3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:297:100
  wire _row_1_d_x2_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:296:100
  wire _row_1_d_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:296:100
  wire _row_1_n_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:295:100
  wire _row_1_n_t2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:294:100
  wire _row_1_d_x1_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:293:100
  wire _row_1_d_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:293:100
  wire _row_1_n_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:292:100
  wire _row_1_n_t1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:291:100
  wire _row_1_d_x0_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:290:100
  wire _row_1_d_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:290:100
  wire _row_1_n_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:289:100
  wire _row_1_d_x8_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:288:100
  wire _row_1_d_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:288:100
  wire _row_1_n_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:287:100
  wire _row_1_d_x7_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:286:100
  wire _row_1_d_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:286:100
  wire _row_1_n_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:285:100
  wire _row_1_n_t7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:284:100
  wire _row_1_d_x6_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:283:100
  wire _row_1_d_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:283:100
  wire _row_1_n_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:282:100
  wire _row_1_n_t6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:281:100
  wire _row_1_d_x8_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:280:100
  wire _row_1_d_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:280:100
  wire _row_1_n_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:279:100
  wire _row_1_n_t8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:278:100
  wire _row_1_d_x5_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:277:100
  wire _row_1_d_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:277:100
  wire _row_1_n_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:276:100
  wire _row_1_n_t5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:275:100
  wire _row_1_d_x4_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:274:100
  wire _row_1_d_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:274:100
  wire _row_1_n_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:273:100
  wire _row_1_n_t4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:272:100
  wire _row_1_d_x8_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:271:100
  wire _row_1_d_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:271:100
  wire _row_1_n_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:270:100
  wire _row_1_n_t8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:269:100
  wire _row_1_d_x7_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:268:100
  wire _row_1_d_x7_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:268:100
  wire _row_1_d_x6_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:267:100
  wire _row_1_d_x6_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:267:100
  wire _row_1_d_x5_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:266:100
  wire _row_1_d_x5_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:266:100
  wire _row_1_d_x4_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:265:100
  wire _row_1_d_x4_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:265:100
  wire _row_1_d_x3_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:264:100
  wire _row_1_d_x3_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:264:100
  wire _row_1_d_x2_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:263:100
  wire _row_1_d_x2_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:263:100
  wire _row_1_d_x1_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:262:100
  wire _row_1_d_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:262:100
  wire _row_1_d_x0_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:261:100
  wire _row_1_d_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:261:100
  wire _row_1_n_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:260:100
  wire _row_1_n_t0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:259:83
  wire _row_1_n_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:258:83
  wire _row_1_n_w2_add_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:257:85
  wire _row_1_n_w2_sub_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:256:85
  wire _row_1_n_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:255:64
  wire _row_1_n_w3_add_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:254:85
  wire _row_1_n_w3_sub_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:253:85
  wire _row_1_n_w3_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:252:64
  wire _row_1_n_w1_add_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:251:85
  wire _row_1_n_w1_sub_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:250:85
  wire _row_1_n_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:249:64
  wire _row_1_n_c181_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:248:76
  wire _row_1_n_c181_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:247:76
  wire _row_1_n_c128_2_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:246:76
  wire _row_1_n_c128_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:245:76
  wire _row_1_n_c128_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:244:76
  wire _row_0_n_shr_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:243:87
  wire _row_0_n_tmp_7_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:242:105
  wire _row_0_n_shr_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:241:87
  wire _row_0_n_tmp_6_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:240:105
  wire _row_0_n_shr_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:239:87
  wire _row_0_n_tmp_5_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:238:105
  wire _row_0_n_shr_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:237:87
  wire _row_0_n_tmp_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:236:105
  wire _row_0_n_shr_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:235:87
  wire _row_0_n_tmp_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:234:105
  wire _row_0_n_shr_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:233:87
  wire _row_0_n_tmp_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:232:105
  wire _row_0_n_shr_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:231:87
  wire _row_0_n_tmp_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:230:105
  wire _row_0_n_shr_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:229:87
  wire _row_0_n_tmp_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:228:105
  wire _row_0_d_x4_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:227:100
  wire _row_0_d_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:227:100
  wire _row_0_n_x4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:226:83
  wire _row_0_n_w4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:225:100
  wire _row_0_n_v4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:224:100
  wire _row_0_n_u4_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:223:100
  wire _row_0_d_x2_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:222:100
  wire _row_0_d_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:222:100
  wire _row_0_n_x2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:221:83
  wire _row_0_n_w2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:220:100
  wire _row_0_n_v2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:219:100
  wire _row_0_n_u2_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:218:100
  wire _row_0_d_x0_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:217:100
  wire _row_0_d_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:217:100
  wire _row_0_n_x0_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:216:100
  wire _row_0_d_x3_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:215:100
  wire _row_0_d_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:215:100
  wire _row_0_n_x3_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:214:100
  wire _row_0_d_x8_4_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:213:100
  wire _row_0_d_x8_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:213:100
  wire _row_0_n_x8_4_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:212:100
  wire _row_0_d_x7_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:211:100
  wire _row_0_d_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:211:100
  wire _row_0_n_x7_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:210:100
  wire _row_0_d_x5_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:209:100
  wire _row_0_d_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:209:100
  wire _row_0_n_x5_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:208:100
  wire _row_0_d_x6_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:207:100
  wire _row_0_d_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:207:100
  wire _row_0_n_x6_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:206:100
  wire _row_0_d_x4_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:205:100
  wire _row_0_d_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:205:100
  wire _row_0_n_x4_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:204:100
  wire _row_0_d_x1_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:203:100
  wire _row_0_d_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:203:100
  wire _row_0_n_x1_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:202:100
  wire _row_0_d_x3_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:201:100
  wire _row_0_d_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:201:100
  wire _row_0_n_x3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:200:100
  wire _row_0_n_t3_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:199:100
  wire _row_0_d_x2_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:198:100
  wire _row_0_d_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:198:100
  wire _row_0_n_x2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:197:100
  wire _row_0_n_t2_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:196:100
  wire _row_0_d_x1_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:195:100
  wire _row_0_d_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:195:100
  wire _row_0_n_x1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:194:100
  wire _row_0_n_t1_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:193:100
  wire _row_0_d_x0_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:192:100
  wire _row_0_d_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:192:100
  wire _row_0_n_x0_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:191:100
  wire _row_0_d_x8_3_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:190:100
  wire _row_0_d_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:190:100
  wire _row_0_n_x8_3_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:189:100
  wire _row_0_d_x7_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:188:100
  wire _row_0_d_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:188:100
  wire _row_0_n_x7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:187:100
  wire _row_0_n_t7_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:186:100
  wire _row_0_d_x6_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:185:100
  wire _row_0_d_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:185:100
  wire _row_0_n_x6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:184:100
  wire _row_0_n_t6_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:183:100
  wire _row_0_d_x8_2_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:182:100
  wire _row_0_d_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:182:100
  wire _row_0_n_x8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:181:100
  wire _row_0_n_t8_2_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:180:100
  wire _row_0_d_x5_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:179:100
  wire _row_0_d_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:179:100
  wire _row_0_n_x5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:178:100
  wire _row_0_n_t5_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:177:100
  wire _row_0_d_x4_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:176:100
  wire _row_0_d_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:176:100
  wire _row_0_n_x4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:175:100
  wire _row_0_n_t4_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:174:100
  wire _row_0_d_x8_1_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:173:100
  wire _row_0_d_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:173:100
  wire _row_0_n_x8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:172:100
  wire _row_0_n_t8_1_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:171:100
  wire _row_0_d_x7_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:170:100
  wire _row_0_d_x7_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:170:100
  wire _row_0_d_x6_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:169:100
  wire _row_0_d_x6_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:169:100
  wire _row_0_d_x5_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:168:100
  wire _row_0_d_x5_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:168:100
  wire _row_0_d_x4_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:167:100
  wire _row_0_d_x4_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:167:100
  wire _row_0_d_x3_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:166:100
  wire _row_0_d_x3_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:166:100
  wire _row_0_d_x2_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:165:100
  wire _row_0_d_x2_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:165:100
  wire _row_0_d_x1_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:164:100
  wire _row_0_d_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:164:100
  wire _row_0_d_x0_0_y;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:163:100
  wire _row_0_d_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:163:100
  wire _row_0_n_x0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:162:100
  wire _row_0_n_t0_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:161:83
  wire _row_0_n_x1_0_z;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:160:83
  wire _row_0_n_w2_add_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:159:85
  wire _row_0_n_w2_sub_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:158:85
  wire _row_0_n_w6_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:157:64
  wire _row_0_n_w3_add_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:156:85
  wire _row_0_n_w3_sub_w5_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:155:85
  wire _row_0_n_w3_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:154:64
  wire _row_0_n_w1_add_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:153:85
  wire _row_0_n_w1_sub_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:152:85
  wire _row_0_n_w7_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:151:64
  wire _row_0_n_c181_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:150:76
  wire _row_0_n_c181_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:149:76
  wire _row_0_n_c128_2_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:148:76
  wire _row_0_n_c128_1_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:147:76
  wire _row_0_n_c128_0_value;	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:146:76

  C128 row_0_n_c128_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:146:76
    .clock (clock),
    .reset (reset),
    .value (_row_0_n_c128_0_value)
  );
  C128 row_0_n_c128_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:147:76
    .clock (clock),
    .reset (reset),
    .value (_row_0_n_c128_1_value)
  );
  C128 row_0_n_c128_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:148:76
    .clock (clock),
    .reset (reset),
    .value (_row_0_n_c128_2_value)
  );
  C181 row_0_n_c181_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:149:76
    .clock (clock),
    .reset (reset),
    .value (_row_0_n_c181_0_value)
  );
  C181 row_0_n_c181_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:150:76
    .clock (clock),
    .reset (reset),
    .value (_row_0_n_c181_1_value)
  );
  W7 row_0_n_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:151:64
    .clock (clock),
    .reset (reset),
    .value (_row_0_n_w7_value)
  );
  W1_sub_W7 row_0_n_w1_sub_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:152:85
    .clock (clock),
    .reset (reset),
    .value (_row_0_n_w1_sub_w7_value)
  );
  W1_add_W7 row_0_n_w1_add_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:153:85
    .clock (clock),
    .reset (reset),
    .value (_row_0_n_w1_add_w7_value)
  );
  W3 row_0_n_w3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:154:64
    .clock (clock),
    .reset (reset),
    .value (_row_0_n_w3_value)
  );
  W3_sub_W5 row_0_n_w3_sub_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:155:85
    .clock (clock),
    .reset (reset),
    .value (_row_0_n_w3_sub_w5_value)
  );
  W3_add_W5 row_0_n_w3_add_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:156:85
    .clock (clock),
    .reset (reset),
    .value (_row_0_n_w3_add_w5_value)
  );
  W6 row_0_n_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:157:64
    .clock (clock),
    .reset (reset),
    .value (_row_0_n_w6_value)
  );
  W2_sub_W6 row_0_n_w2_sub_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:158:85
    .clock (clock),
    .reset (reset),
    .value (_row_0_n_w2_sub_w6_value)
  );
  W2_add_W6 row_0_n_w2_add_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:159:85
    .clock (clock),
    .reset (reset),
    .value (_row_0_n_w2_add_w6_value)
  );
  SHL_11 row_0_n_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:160:83
    .clock (clock),
    .reset (reset),
    .x     (n_in_0_4_x),
    .z     (_row_0_n_x1_0_z)
  );
  SHL_11 row_0_n_t0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:161:83
    .clock (clock),
    .reset (reset),
    .x     (n_in_0_0_x),
    .z     (_row_0_n_t0_0_z)
  );
  ADD row_0_n_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:162:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_t0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:161:83
    .y     (_row_0_n_c128_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:146:76
    .z     (_row_0_n_x0_0_z)
  );
  dup_2 row_0_d_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:163:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:162:100
    .y     (_row_0_d_x0_0_y),
    .z     (_row_0_d_x0_0_z)
  );
  dup_2 row_0_d_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:164:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:160:83
    .y     (_row_0_d_x1_0_y),
    .z     (_row_0_d_x1_0_z)
  );
  dup_2 row_0_d_x2_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:165:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_0_6_x),
    .y     (_row_0_d_x2_0_y),
    .z     (_row_0_d_x2_0_z)
  );
  dup_2 row_0_d_x3_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:166:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_0_2_x),
    .y     (_row_0_d_x3_0_y),
    .z     (_row_0_d_x3_0_z)
  );
  dup_2 row_0_d_x4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:167:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_0_1_x),
    .y     (_row_0_d_x4_0_y),
    .z     (_row_0_d_x4_0_z)
  );
  dup_2 row_0_d_x5_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:168:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_0_7_x),
    .y     (_row_0_d_x5_0_y),
    .z     (_row_0_d_x5_0_z)
  );
  dup_2 row_0_d_x6_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:169:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_0_5_x),
    .y     (_row_0_d_x6_0_y),
    .z     (_row_0_d_x6_0_z)
  );
  dup_2 row_0_d_x7_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:170:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_0_3_x),
    .y     (_row_0_d_x7_0_y),
    .z     (_row_0_d_x7_0_z)
  );
  ADD row_0_n_t8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:171:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_45_2295_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2313:114
    .y     (_row_0_d_x5_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:168:100
    .z     (_row_0_n_t8_1_z)
  );
  MUL row_0_n_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:172:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:151:64
    .y     (_row_0_n_t8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:171:100
    .z     (_row_0_n_x8_1_z)
  );
  dup_2 row_0_d_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:173:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:172:100
    .y     (_row_0_d_x8_1_y),
    .z     (_row_0_d_x8_1_z)
  );
  MUL row_0_n_t4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:174:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_w1_sub_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:152:85
    .y     (_row_0_d_x4_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:167:100
    .z     (_row_0_n_t4_1_z)
  );
  ADD row_0_n_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:175:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x8_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:173:100
    .y     (_delay_INT16_200_2293_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2311:118
    .z     (_row_0_n_x4_1_z)
  );
  dup_2 row_0_d_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:176:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:175:100
    .y     (_row_0_d_x4_1_y),
    .z     (_row_0_d_x4_1_z)
  );
  MUL row_0_n_t5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:177:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_w1_add_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:153:85
    .y     (_row_0_d_x5_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:168:100
    .z     (_row_0_n_t5_1_z)
  );
  SUB row_0_n_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:178:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:173:100
    .y     (_delay_INT16_149_2292_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2310:118
    .z     (_row_0_n_x5_1_z)
  );
  dup_2 row_0_d_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:179:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:178:100
    .y     (_row_0_d_x5_1_y),
    .z     (_row_0_d_x5_1_z)
  );
  ADD row_0_n_t8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:180:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x6_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:169:100
    .y     (_delay_INT16_24_2291_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2309:114
    .z     (_row_0_n_t8_2_z)
  );
  MUL row_0_n_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:181:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_w3_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:154:64
    .y     (_row_0_n_t8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:180:100
    .z     (_row_0_n_x8_2_z)
  );
  dup_2 row_0_d_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:182:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:181:100
    .y     (_row_0_d_x8_2_y),
    .z     (_row_0_d_x8_2_z)
  );
  MUL row_0_n_t6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:183:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_w3_sub_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:155:85
    .y     (_row_0_d_x6_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:169:100
    .z     (_row_0_n_t6_1_z)
  );
  SUB row_0_n_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:184:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x8_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:182:100
    .y     (_delay_INT16_171_2290_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2308:118
    .z     (_row_0_n_x6_1_z)
  );
  dup_2 row_0_d_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:185:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:184:100
    .y     (_row_0_d_x6_1_y),
    .z     (_row_0_d_x6_1_z)
  );
  MUL row_0_n_t7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:186:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_w3_add_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:156:85
    .y     (_delay_INT16_15_2289_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2307:114
    .z     (_row_0_n_t7_1_z)
  );
  SUB row_0_n_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:187:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:182:100
    .y     (_delay_INT16_93_2288_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2306:114
    .z     (_row_0_n_x7_1_z)
  );
  dup_2 row_0_d_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:188:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:187:100
    .y     (_row_0_d_x7_1_y),
    .z     (_row_0_d_x7_1_z)
  );
  ADD row_0_n_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:189:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x0_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:163:100
    .y     (_delay_INT16_29_2301_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2319:114
    .z     (_row_0_n_x8_3_z)
  );
  dup_2 row_0_d_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:190:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:189:100
    .y     (_row_0_d_x8_3_y),
    .z     (_row_0_d_x8_3_z)
  );
  SUB row_0_n_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:191:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:163:100
    .y     (_delay_INT16_29_2287_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2305:114
    .z     (_row_0_n_x0_1_z)
  );
  dup_2 row_0_d_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:192:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:191:100
    .y     (_row_0_d_x0_1_y),
    .z     (_row_0_d_x0_1_z)
  );
  ADD row_0_n_t1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:193:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x3_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:166:100
    .y     (_delay_INT16_100_2285_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2303:118
    .z     (_row_0_n_t1_1_z)
  );
  MUL row_0_n_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:194:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:157:64
    .y     (_row_0_n_t1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:193:100
    .z     (_row_0_n_x1_1_z)
  );
  dup_2 row_0_d_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:195:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:194:100
    .y     (_row_0_d_x1_1_y),
    .z     (_row_0_d_x1_1_z)
  );
  MUL row_0_n_t2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:196:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_w2_add_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:159:85
    .y     (_delay_INT16_27_2283_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2301:114
    .z     (_row_0_n_t2_1_z)
  );
  SUB row_0_n_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:197:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x1_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:195:100
    .y     (_delay_INT16_147_2282_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2300:118
    .z     (_row_0_n_x2_1_z)
  );
  dup_2 row_0_d_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:198:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:197:100
    .y     (_row_0_d_x2_1_y),
    .z     (_row_0_d_x2_1_z)
  );
  MUL row_0_n_t3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:199:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_w2_sub_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:158:85
    .y     (_row_0_d_x3_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:166:100
    .z     (_row_0_n_t3_1_z)
  );
  ADD row_0_n_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:200:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:195:100
    .y     (_delay_INT16_127_2281_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2299:118
    .z     (_row_0_n_x3_1_z)
  );
  dup_2 row_0_d_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:201:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:200:100
    .y     (_row_0_d_x3_1_y),
    .z     (_row_0_d_x3_1_z)
  );
  ADD row_0_n_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:202:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x4_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:176:100
    .y     (_delay_INT16_42_2279_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2297:114
    .z     (_row_0_n_x1_2_z)
  );
  dup_2 row_0_d_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:203:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:202:100
    .y     (_row_0_d_x1_2_y),
    .z     (_row_0_d_x1_2_z)
  );
  SUB row_0_n_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:204:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:176:100
    .y     (_delay_INT16_42_2277_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2295:114
    .z     (_row_0_n_x4_2_z)
  );
  dup_2 row_0_d_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:205:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:204:100
    .y     (_row_0_d_x4_2_y),
    .z     (_row_0_d_x4_2_z)
  );
  ADD row_0_n_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:206:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x5_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:179:100
    .y     (_delay_INT16_65_2276_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2294:114
    .z     (_row_0_n_x6_2_z)
  );
  dup_2 row_0_d_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:207:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:206:100
    .y     (_row_0_d_x6_2_y),
    .z     (_row_0_d_x6_2_z)
  );
  SUB row_0_n_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:208:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:179:100
    .y     (_delay_INT16_65_2275_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2293:114
    .z     (_row_0_n_x5_2_z)
  );
  dup_2 row_0_d_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:209:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:208:100
    .y     (_row_0_d_x5_2_y),
    .z     (_row_0_d_x5_2_z)
  );
  ADD row_0_n_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:210:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_162_2274_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2292:118
    .y     (_row_0_d_x3_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:201:100
    .z     (_row_0_n_x7_2_z)
  );
  dup_2 row_0_d_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:211:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:210:100
    .y     (_row_0_d_x7_2_y),
    .z     (_row_0_d_x7_2_z)
  );
  SUB row_0_n_x8_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:212:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_162_2273_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2291:118
    .y     (_row_0_d_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:201:100
    .z     (_row_0_n_x8_4_z)
  );
  dup_2 row_0_d_x8_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:213:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x8_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:212:100
    .y     (_row_0_d_x8_4_y),
    .z     (_row_0_d_x8_4_z)
  );
  ADD row_0_n_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:214:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_106_2297_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2315:118
    .y     (_row_0_d_x2_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:198:100
    .z     (_row_0_n_x3_2_z)
  );
  dup_2 row_0_d_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:215:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:214:100
    .y     (_row_0_d_x3_2_y),
    .z     (_row_0_d_x3_2_z)
  );
  SUB row_0_n_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:216:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_106_2271_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2289:118
    .y     (_row_0_d_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:198:100
    .z     (_row_0_n_x0_2_z)
  );
  dup_2 row_0_d_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:217:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:216:100
    .y     (_row_0_d_x0_2_y),
    .z     (_row_0_d_x0_2_z)
  );
  ADD row_0_n_u2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:218:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_89_2270_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2288:114
    .y     (_row_0_d_x5_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:209:100
    .z     (_row_0_n_u2_2_z)
  );
  MUL row_0_n_v2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:219:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_c181_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:149:76
    .y     (_row_0_n_u2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:218:100
    .z     (_row_0_n_v2_2_z)
  );
  ADD row_0_n_w2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:220:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_v2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:219:100
    .y     (_row_0_n_c128_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:147:76
    .z     (_row_0_n_w2_2_z)
  );
  SHR_8 row_0_n_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:221:83
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_w2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:220:100
    .z     (_row_0_n_x2_2_z)
  );
  dup_2 row_0_d_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:222:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:221:83
    .y     (_row_0_d_x2_2_y),
    .z     (_row_0_d_x2_2_z)
  );
  SUB row_0_n_u4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:223:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_89_2269_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2287:114
    .y     (_row_0_d_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:209:100
    .z     (_row_0_n_u4_3_z)
  );
  MUL row_0_n_v4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:224:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_c181_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:150:76
    .y     (_row_0_n_u4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:223:100
    .z     (_row_0_n_v4_3_z)
  );
  ADD row_0_n_w4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:225:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_v4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:224:100
    .y     (_row_0_n_c128_2_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:148:76
    .z     (_row_0_n_w4_3_z)
  );
  SHR_8 row_0_n_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:226:83
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_w4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:225:100
    .z     (_row_0_n_x4_3_z)
  );
  dup_2 row_0_d_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:227:100
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:226:83
    .y     (_row_0_d_x4_3_y),
    .z     (_row_0_d_x4_3_z)
  );
  ADD row_0_n_tmp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:228:105
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x7_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:211:100
    .y     (_delay_INT16_20_2267_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2285:114
    .z     (_row_0_n_tmp_0_z)
  );
  SHR_8 row_0_n_shr_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:229:87
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_tmp_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:228:105
    .z     (_row_0_n_shr_0_z)
  );
  ADD row_0_n_tmp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:230:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_206_2266_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2284:118
    .y     (_row_0_d_x2_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:222:100
    .z     (_row_0_n_tmp_1_z)
  );
  SHR_8 row_0_n_shr_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:231:87
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_tmp_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:230:105
    .z     (_row_0_n_shr_1_z)
  );
  ADD row_0_n_tmp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:232:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_162_2264_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2282:118
    .y     (_row_0_d_x4_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:227:100
    .z     (_row_0_n_tmp_2_z)
  );
  SHR_8 row_0_n_shr_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:233:87
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_tmp_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:232:105
    .z     (_row_0_n_shr_2_z)
  );
  ADD row_0_n_tmp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:234:105
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x8_4_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:213:100
    .y     (_delay_INT16_49_2263_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2281:114
    .z     (_row_0_n_tmp_3_z)
  );
  SHR_8 row_0_n_shr_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:235:87
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_tmp_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:234:105
    .z     (_row_0_n_shr_3_z)
  );
  SUB row_0_n_tmp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:236:105
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x8_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:213:100
    .y     (_delay_INT16_49_2323_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2341:114
    .z     (_row_0_n_tmp_4_z)
  );
  SHR_8 row_0_n_shr_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:237:87
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_tmp_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:236:105
    .z     (_row_0_n_shr_4_z)
  );
  SUB row_0_n_tmp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:238:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_162_2262_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2280:118
    .y     (_row_0_d_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:227:100
    .z     (_row_0_n_tmp_5_z)
  );
  SHR_8 row_0_n_shr_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:239:87
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_tmp_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:238:105
    .z     (_row_0_n_shr_5_z)
  );
  SUB row_0_n_tmp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:240:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_206_2261_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2279:118
    .y     (_row_0_d_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:222:100
    .z     (_row_0_n_tmp_6_z)
  );
  SHR_8 row_0_n_shr_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:241:87
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_tmp_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:240:105
    .z     (_row_0_n_shr_6_z)
  );
  SUB row_0_n_tmp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:242:105
    .clock (clock),
    .reset (reset),
    .x     (_row_0_d_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:211:100
    .y     (_delay_INT16_20_2260_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2278:114
    .z     (_row_0_n_tmp_7_z)
  );
  SHR_8 row_0_n_shr_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:243:87
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_tmp_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:242:105
    .z     (_row_0_n_shr_7_z)
  );
  C128 row_1_n_c128_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:244:76
    .clock (clock),
    .reset (reset),
    .value (_row_1_n_c128_0_value)
  );
  C128 row_1_n_c128_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:245:76
    .clock (clock),
    .reset (reset),
    .value (_row_1_n_c128_1_value)
  );
  C128 row_1_n_c128_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:246:76
    .clock (clock),
    .reset (reset),
    .value (_row_1_n_c128_2_value)
  );
  C181 row_1_n_c181_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:247:76
    .clock (clock),
    .reset (reset),
    .value (_row_1_n_c181_0_value)
  );
  C181 row_1_n_c181_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:248:76
    .clock (clock),
    .reset (reset),
    .value (_row_1_n_c181_1_value)
  );
  W7 row_1_n_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:249:64
    .clock (clock),
    .reset (reset),
    .value (_row_1_n_w7_value)
  );
  W1_sub_W7 row_1_n_w1_sub_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:250:85
    .clock (clock),
    .reset (reset),
    .value (_row_1_n_w1_sub_w7_value)
  );
  W1_add_W7 row_1_n_w1_add_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:251:85
    .clock (clock),
    .reset (reset),
    .value (_row_1_n_w1_add_w7_value)
  );
  W3 row_1_n_w3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:252:64
    .clock (clock),
    .reset (reset),
    .value (_row_1_n_w3_value)
  );
  W3_sub_W5 row_1_n_w3_sub_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:253:85
    .clock (clock),
    .reset (reset),
    .value (_row_1_n_w3_sub_w5_value)
  );
  W3_add_W5 row_1_n_w3_add_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:254:85
    .clock (clock),
    .reset (reset),
    .value (_row_1_n_w3_add_w5_value)
  );
  W6 row_1_n_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:255:64
    .clock (clock),
    .reset (reset),
    .value (_row_1_n_w6_value)
  );
  W2_sub_W6 row_1_n_w2_sub_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:256:85
    .clock (clock),
    .reset (reset),
    .value (_row_1_n_w2_sub_w6_value)
  );
  W2_add_W6 row_1_n_w2_add_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:257:85
    .clock (clock),
    .reset (reset),
    .value (_row_1_n_w2_add_w6_value)
  );
  SHL_11 row_1_n_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:258:83
    .clock (clock),
    .reset (reset),
    .x     (n_in_1_4_x),
    .z     (_row_1_n_x1_0_z)
  );
  SHL_11 row_1_n_t0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:259:83
    .clock (clock),
    .reset (reset),
    .x     (n_in_1_0_x),
    .z     (_row_1_n_t0_0_z)
  );
  ADD row_1_n_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:260:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_t0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:259:83
    .y     (_row_1_n_c128_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:244:76
    .z     (_row_1_n_x0_0_z)
  );
  dup_2 row_1_d_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:261:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:260:100
    .y     (_row_1_d_x0_0_y),
    .z     (_row_1_d_x0_0_z)
  );
  dup_2 row_1_d_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:262:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:258:83
    .y     (_row_1_d_x1_0_y),
    .z     (_row_1_d_x1_0_z)
  );
  dup_2 row_1_d_x2_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:263:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_1_6_x),
    .y     (_row_1_d_x2_0_y),
    .z     (_row_1_d_x2_0_z)
  );
  dup_2 row_1_d_x3_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:264:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_1_2_x),
    .y     (_row_1_d_x3_0_y),
    .z     (_row_1_d_x3_0_z)
  );
  dup_2 row_1_d_x4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:265:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_1_1_x),
    .y     (_row_1_d_x4_0_y),
    .z     (_row_1_d_x4_0_z)
  );
  dup_2 row_1_d_x5_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:266:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_1_7_x),
    .y     (_row_1_d_x5_0_y),
    .z     (_row_1_d_x5_0_z)
  );
  dup_2 row_1_d_x6_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:267:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_1_5_x),
    .y     (_row_1_d_x6_0_y),
    .z     (_row_1_d_x6_0_z)
  );
  dup_2 row_1_d_x7_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:268:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_1_3_x),
    .y     (_row_1_d_x7_0_y),
    .z     (_row_1_d_x7_0_z)
  );
  ADD row_1_n_t8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:269:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_d_x4_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:265:100
    .y     (_delay_INT16_23_2257_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2275:114
    .z     (_row_1_n_t8_1_z)
  );
  MUL row_1_n_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:270:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:249:64
    .y     (_row_1_n_t8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:269:100
    .z     (_row_1_n_x8_1_z)
  );
  dup_2 row_1_d_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:271:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:270:100
    .y     (_row_1_d_x8_1_y),
    .z     (_row_1_d_x8_1_z)
  );
  MUL row_1_n_t4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:272:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_w1_sub_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:250:85
    .y     (_row_1_d_x4_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:265:100
    .z     (_row_1_n_t4_1_z)
  );
  ADD row_1_n_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:273:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_d_x8_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:271:100
    .y     (_delay_INT16_26_2256_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2274:114
    .z     (_row_1_n_x4_1_z)
  );
  dup_2 row_1_d_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:274:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:273:100
    .y     (_row_1_d_x4_1_y),
    .z     (_row_1_d_x4_1_z)
  );
  MUL row_1_n_t5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:275:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_w1_add_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:251:85
    .y     (_row_1_d_x5_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:266:100
    .z     (_row_1_n_t5_1_z)
  );
  SUB row_1_n_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:276:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_d_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:271:100
    .y     (_delay_INT16_97_2255_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2273:114
    .z     (_row_1_n_x5_1_z)
  );
  dup_2 row_1_d_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:277:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:276:100
    .y     (_row_1_d_x5_1_y),
    .z     (_row_1_d_x5_1_z)
  );
  ADD row_1_n_t8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:278:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_29_2253_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2271:114
    .y     (_row_1_d_x7_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:268:100
    .z     (_row_1_n_t8_2_z)
  );
  MUL row_1_n_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:279:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_w3_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:252:64
    .y     (_row_1_n_t8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:278:100
    .z     (_row_1_n_x8_2_z)
  );
  dup_2 row_1_d_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:280:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:279:100
    .y     (_row_1_d_x8_2_y),
    .z     (_row_1_d_x8_2_z)
  );
  MUL row_1_n_t6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:281:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_w3_sub_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:253:85
    .y     (_row_1_d_x6_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:267:100
    .z     (_row_1_n_t6_1_z)
  );
  SUB row_1_n_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:282:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_d_x8_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:280:100
    .y     (_delay_INT16_109_2252_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2270:118
    .z     (_row_1_n_x6_1_z)
  );
  dup_2 row_1_d_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:283:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:282:100
    .y     (_row_1_d_x6_1_y),
    .z     (_row_1_d_x6_1_z)
  );
  MUL row_1_n_t7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:284:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_w3_add_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:254:85
    .y     (_row_1_d_x7_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:268:100
    .z     (_row_1_n_t7_1_z)
  );
  SUB row_1_n_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:285:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_d_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:280:100
    .y     (_delay_INT16_89_2250_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2268:114
    .z     (_row_1_n_x7_1_z)
  );
  dup_2 row_1_d_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:286:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:285:100
    .y     (_row_1_d_x7_1_y),
    .z     (_row_1_d_x7_1_z)
  );
  ADD row_1_n_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:287:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_d_x0_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:261:100
    .y     (_delay_INT16_61_2249_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2267:114
    .z     (_row_1_n_x8_3_z)
  );
  dup_2 row_1_d_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:288:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:287:100
    .y     (_row_1_d_x8_3_y),
    .z     (_row_1_d_x8_3_z)
  );
  SUB row_1_n_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:289:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_d_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:261:100
    .y     (_delay_INT16_61_2247_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2265:114
    .z     (_row_1_n_x0_1_z)
  );
  dup_2 row_1_d_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:290:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:289:100
    .y     (_row_1_d_x0_1_y),
    .z     (_row_1_d_x0_1_z)
  );
  ADD row_1_n_t1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:291:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_d_x3_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:264:100
    .y     (_delay_INT16_10_2246_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2264:114
    .z     (_row_1_n_t1_1_z)
  );
  MUL row_1_n_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:292:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:255:64
    .y     (_row_1_n_t1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:291:100
    .z     (_row_1_n_x1_1_z)
  );
  dup_2 row_1_d_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:293:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:292:100
    .y     (_row_1_d_x1_1_y),
    .z     (_row_1_d_x1_1_z)
  );
  MUL row_1_n_t2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:294:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_w2_add_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:257:85
    .y     (_row_1_d_x2_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:263:100
    .z     (_row_1_n_t2_1_z)
  );
  SUB row_1_n_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:295:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_d_x1_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:293:100
    .y     (_delay_INT16_139_2245_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2263:118
    .z     (_row_1_n_x2_1_z)
  );
  dup_2 row_1_d_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:296:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:295:100
    .y     (_row_1_d_x2_1_y),
    .z     (_row_1_d_x2_1_z)
  );
  MUL row_1_n_t3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:297:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_w2_sub_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:256:85
    .y     (_row_1_d_x3_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:264:100
    .z     (_row_1_n_t3_1_z)
  );
  ADD row_1_n_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:298:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_d_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:293:100
    .y     (_delay_INT16_61_2244_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2262:114
    .z     (_row_1_n_x3_1_z)
  );
  dup_2 row_1_d_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:299:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:298:100
    .y     (_row_1_d_x3_1_y),
    .z     (_row_1_d_x3_1_z)
  );
  ADD row_1_n_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:300:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_85_2243_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2261:114
    .y     (_row_1_d_x6_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:283:100
    .z     (_row_1_n_x1_2_z)
  );
  dup_2 row_1_d_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:301:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:300:100
    .y     (_row_1_d_x1_2_y),
    .z     (_row_1_d_x1_2_z)
  );
  SUB row_1_n_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:302:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_85_2242_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2260:114
    .y     (_row_1_d_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:283:100
    .z     (_row_1_n_x4_2_z)
  );
  dup_2 row_1_d_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:303:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:302:100
    .y     (_row_1_d_x4_2_y),
    .z     (_row_1_d_x4_2_z)
  );
  ADD row_1_n_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:304:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_126_2241_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2259:118
    .y     (_row_1_d_x7_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:286:100
    .z     (_row_1_n_x6_2_z)
  );
  dup_2 row_1_d_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:305:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:304:100
    .y     (_row_1_d_x6_2_y),
    .z     (_row_1_d_x6_2_z)
  );
  SUB row_1_n_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:306:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_126_2240_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2258:118
    .y     (_row_1_d_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:286:100
    .z     (_row_1_n_x5_2_z)
  );
  dup_2 row_1_d_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:307:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:306:100
    .y     (_row_1_d_x5_2_y),
    .z     (_row_1_d_x5_2_z)
  );
  ADD row_1_n_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:308:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_85_2239_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2257:114
    .y     (_row_1_d_x3_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:299:100
    .z     (_row_1_n_x7_2_z)
  );
  dup_2 row_1_d_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:309:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:308:100
    .y     (_row_1_d_x7_2_y),
    .z     (_row_1_d_x7_2_z)
  );
  SUB row_1_n_x8_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:310:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_85_2238_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2256:114
    .y     (_row_1_d_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:299:100
    .z     (_row_1_n_x8_4_z)
  );
  dup_2 row_1_d_x8_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:311:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x8_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:310:100
    .y     (_row_1_d_x8_4_y),
    .z     (_row_1_d_x8_4_z)
  );
  ADD row_1_n_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:312:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_153_2237_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2255:118
    .y     (_row_1_d_x2_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:296:100
    .z     (_row_1_n_x3_2_z)
  );
  dup_2 row_1_d_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:313:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:312:100
    .y     (_row_1_d_x3_2_y),
    .z     (_row_1_d_x3_2_z)
  );
  SUB row_1_n_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:314:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_153_2236_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2254:118
    .y     (_row_1_d_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:296:100
    .z     (_row_1_n_x0_2_z)
  );
  dup_2 row_1_d_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:315:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:314:100
    .y     (_row_1_d_x0_2_y),
    .z     (_row_1_d_x0_2_z)
  );
  ADD row_1_n_u2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:316:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_48_2234_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2252:114
    .y     (_row_1_d_x5_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:307:100
    .z     (_row_1_n_u2_2_z)
  );
  MUL row_1_n_v2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:317:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_c181_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:247:76
    .y     (_row_1_n_u2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:316:100
    .z     (_row_1_n_v2_2_z)
  );
  ADD row_1_n_w2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:318:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_v2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:317:100
    .y     (_row_1_n_c128_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:245:76
    .z     (_row_1_n_w2_2_z)
  );
  SHR_8 row_1_n_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:319:83
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_w2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:318:100
    .z     (_row_1_n_x2_2_z)
  );
  dup_2 row_1_d_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:320:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:319:83
    .y     (_row_1_d_x2_2_y),
    .z     (_row_1_d_x2_2_z)
  );
  SUB row_1_n_u4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:321:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_48_2233_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2251:114
    .y     (_row_1_d_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:307:100
    .z     (_row_1_n_u4_3_z)
  );
  MUL row_1_n_v4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:322:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_c181_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:248:76
    .y     (_row_1_n_u4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:321:100
    .z     (_row_1_n_v4_3_z)
  );
  ADD row_1_n_w4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:323:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_v4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:322:100
    .y     (_row_1_n_c128_2_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:246:76
    .z     (_row_1_n_w4_3_z)
  );
  SHR_8 row_1_n_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:324:83
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_w4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:323:100
    .z     (_row_1_n_x4_3_z)
  );
  dup_2 row_1_d_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:325:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:324:83
    .y     (_row_1_d_x4_3_y),
    .z     (_row_1_d_x4_3_z)
  );
  ADD row_1_n_tmp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:326:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_18_2229_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2247:114
    .y     (_row_1_d_x1_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:301:100
    .z     (_row_1_n_tmp_0_z)
  );
  SHR_8 row_1_n_shr_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:327:87
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_tmp_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:326:105
    .z     (_row_1_n_shr_0_z)
  );
  ADD row_1_n_tmp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:328:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_268_2228_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2246:118
    .y     (_row_1_d_x2_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:320:100
    .z     (_row_1_n_tmp_1_z)
  );
  SHR_8 row_1_n_shr_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:329:87
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_tmp_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:328:105
    .z     (_row_1_n_shr_1_z)
  );
  ADD row_1_n_tmp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:330:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_303_2227_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2245:118
    .y     (_row_1_d_x4_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:325:100
    .z     (_row_1_n_tmp_2_z)
  );
  SHR_8 row_1_n_shr_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:331:87
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_tmp_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:330:105
    .z     (_row_1_n_shr_2_z)
  );
  ADD row_1_n_tmp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:332:105
    .clock (clock),
    .reset (reset),
    .x     (_row_1_d_x8_4_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:311:100
    .y     (_delay_INT16_70_2226_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2244:114
    .z     (_row_1_n_tmp_3_z)
  );
  SHR_8 row_1_n_shr_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:333:87
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_tmp_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:332:105
    .z     (_row_1_n_shr_3_z)
  );
  SUB row_1_n_tmp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:334:105
    .clock (clock),
    .reset (reset),
    .x     (_row_1_d_x8_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:311:100
    .y     (_delay_INT16_70_2235_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2253:114
    .z     (_row_1_n_tmp_4_z)
  );
  SHR_8 row_1_n_shr_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:335:87
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_tmp_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:334:105
    .z     (_row_1_n_shr_4_z)
  );
  SUB row_1_n_tmp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:336:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_303_2222_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2240:118
    .y     (_row_1_d_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:325:100
    .z     (_row_1_n_tmp_5_z)
  );
  SHR_8 row_1_n_shr_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:337:87
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_tmp_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:336:105
    .z     (_row_1_n_shr_5_z)
  );
  SUB row_1_n_tmp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:338:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_268_2221_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2239:118
    .y     (_row_1_d_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:320:100
    .z     (_row_1_n_tmp_6_z)
  );
  SHR_8 row_1_n_shr_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:339:87
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_tmp_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:338:105
    .z     (_row_1_n_shr_6_z)
  );
  SUB row_1_n_tmp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:340:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_18_2219_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2237:114
    .y     (_row_1_d_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:301:100
    .z     (_row_1_n_tmp_7_z)
  );
  SHR_8 row_1_n_shr_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:341:87
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_tmp_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:340:105
    .z     (_row_1_n_shr_7_z)
  );
  C128 row_2_n_c128_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:342:76
    .clock (clock),
    .reset (reset),
    .value (_row_2_n_c128_0_value)
  );
  C128 row_2_n_c128_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:343:76
    .clock (clock),
    .reset (reset),
    .value (_row_2_n_c128_1_value)
  );
  C128 row_2_n_c128_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:344:76
    .clock (clock),
    .reset (reset),
    .value (_row_2_n_c128_2_value)
  );
  C181 row_2_n_c181_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:345:76
    .clock (clock),
    .reset (reset),
    .value (_row_2_n_c181_0_value)
  );
  C181 row_2_n_c181_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:346:76
    .clock (clock),
    .reset (reset),
    .value (_row_2_n_c181_1_value)
  );
  W7 row_2_n_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:347:64
    .clock (clock),
    .reset (reset),
    .value (_row_2_n_w7_value)
  );
  W1_sub_W7 row_2_n_w1_sub_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:348:85
    .clock (clock),
    .reset (reset),
    .value (_row_2_n_w1_sub_w7_value)
  );
  W1_add_W7 row_2_n_w1_add_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:349:85
    .clock (clock),
    .reset (reset),
    .value (_row_2_n_w1_add_w7_value)
  );
  W3 row_2_n_w3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:350:64
    .clock (clock),
    .reset (reset),
    .value (_row_2_n_w3_value)
  );
  W3_sub_W5 row_2_n_w3_sub_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:351:85
    .clock (clock),
    .reset (reset),
    .value (_row_2_n_w3_sub_w5_value)
  );
  W3_add_W5 row_2_n_w3_add_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:352:85
    .clock (clock),
    .reset (reset),
    .value (_row_2_n_w3_add_w5_value)
  );
  W6 row_2_n_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:353:64
    .clock (clock),
    .reset (reset),
    .value (_row_2_n_w6_value)
  );
  W2_sub_W6 row_2_n_w2_sub_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:354:85
    .clock (clock),
    .reset (reset),
    .value (_row_2_n_w2_sub_w6_value)
  );
  W2_add_W6 row_2_n_w2_add_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:355:85
    .clock (clock),
    .reset (reset),
    .value (_row_2_n_w2_add_w6_value)
  );
  SHL_11 row_2_n_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:356:83
    .clock (clock),
    .reset (reset),
    .x     (n_in_2_4_x),
    .z     (_row_2_n_x1_0_z)
  );
  SHL_11 row_2_n_t0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:357:83
    .clock (clock),
    .reset (reset),
    .x     (n_in_2_0_x),
    .z     (_row_2_n_t0_0_z)
  );
  ADD row_2_n_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:358:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_t0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:357:83
    .y     (_row_2_n_c128_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:342:76
    .z     (_row_2_n_x0_0_z)
  );
  dup_2 row_2_d_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:359:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:358:100
    .y     (_row_2_d_x0_0_y),
    .z     (_row_2_d_x0_0_z)
  );
  dup_2 row_2_d_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:360:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:356:83
    .y     (_row_2_d_x1_0_y),
    .z     (_row_2_d_x1_0_z)
  );
  dup_2 row_2_d_x2_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:361:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_2_6_x),
    .y     (_row_2_d_x2_0_y),
    .z     (_row_2_d_x2_0_z)
  );
  dup_2 row_2_d_x3_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:362:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_2_2_x),
    .y     (_row_2_d_x3_0_y),
    .z     (_row_2_d_x3_0_z)
  );
  dup_2 row_2_d_x4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:363:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_2_1_x),
    .y     (_row_2_d_x4_0_y),
    .z     (_row_2_d_x4_0_z)
  );
  dup_2 row_2_d_x5_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:364:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_2_7_x),
    .y     (_row_2_d_x5_0_y),
    .z     (_row_2_d_x5_0_z)
  );
  dup_2 row_2_d_x6_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:365:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_2_5_x),
    .y     (_row_2_d_x6_0_y),
    .z     (_row_2_d_x6_0_z)
  );
  dup_2 row_2_d_x7_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:366:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_2_3_x),
    .y     (_row_2_d_x7_0_y),
    .z     (_row_2_d_x7_0_z)
  );
  ADD row_2_n_t8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:367:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_d_x4_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:363:100
    .y     (_delay_INT16_36_2215_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2233:114
    .z     (_row_2_n_t8_1_z)
  );
  MUL row_2_n_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:368:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:347:64
    .y     (_row_2_n_t8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:367:100
    .z     (_row_2_n_x8_1_z)
  );
  dup_2 row_2_d_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:369:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:368:100
    .y     (_row_2_d_x8_1_y),
    .z     (_row_2_d_x8_1_z)
  );
  MUL row_2_n_t4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:370:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_w1_sub_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:348:85
    .y     (_row_2_d_x4_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:363:100
    .z     (_row_2_n_t4_1_z)
  );
  ADD row_2_n_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:371:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_d_x8_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:369:100
    .y     (_delay_INT16_10_2214_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2232:114
    .z     (_row_2_n_x4_1_z)
  );
  dup_2 row_2_d_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:372:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:371:100
    .y     (_row_2_d_x4_1_y),
    .z     (_row_2_d_x4_1_z)
  );
  MUL row_2_n_t5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:373:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_w1_add_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:349:85
    .y     (_row_2_d_x5_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:364:100
    .z     (_row_2_n_t5_1_z)
  );
  SUB row_2_n_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:374:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_d_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:369:100
    .y     (_delay_INT16_104_2303_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2321:118
    .z     (_row_2_n_x5_1_z)
  );
  dup_2 row_2_d_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:375:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:374:100
    .y     (_row_2_d_x5_1_y),
    .z     (_row_2_d_x5_1_z)
  );
  ADD row_2_n_t8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:376:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_7_2296_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2314:110
    .y     (_row_2_d_x7_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:366:100
    .z     (_row_2_n_t8_2_z)
  );
  MUL row_2_n_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:377:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_w3_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:350:64
    .y     (_row_2_n_t8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:376:100
    .z     (_row_2_n_x8_2_z)
  );
  dup_2 row_2_d_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:378:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:377:100
    .y     (_row_2_d_x8_2_y),
    .z     (_row_2_d_x8_2_z)
  );
  MUL row_2_n_t6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:379:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_w3_sub_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:351:85
    .y     (_row_2_d_x6_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:365:100
    .z     (_row_2_n_t6_1_z)
  );
  SUB row_2_n_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:380:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_d_x8_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:378:100
    .y     (_delay_INT16_149_2213_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2231:118
    .z     (_row_2_n_x6_1_z)
  );
  dup_2 row_2_d_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:381:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:380:100
    .y     (_row_2_d_x6_1_y),
    .z     (_row_2_d_x6_1_z)
  );
  MUL row_2_n_t7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:382:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_w3_add_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:352:85
    .y     (_row_2_d_x7_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:366:100
    .z     (_row_2_n_t7_1_z)
  );
  SUB row_2_n_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:383:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_d_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:378:100
    .y     (_delay_INT16_161_2211_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2229:118
    .z     (_row_2_n_x7_1_z)
  );
  dup_2 row_2_d_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:384:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:383:100
    .y     (_row_2_d_x7_1_y),
    .z     (_row_2_d_x7_1_z)
  );
  ADD row_2_n_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:385:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_117_2210_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2228:118
    .y     (_row_2_d_x1_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:360:100
    .z     (_row_2_n_x8_3_z)
  );
  dup_2 row_2_d_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:386:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:385:100
    .y     (_row_2_d_x8_3_y),
    .z     (_row_2_d_x8_3_z)
  );
  SUB row_2_n_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:387:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_117_2208_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2226:118
    .y     (_row_2_d_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:360:100
    .z     (_row_2_n_x0_1_z)
  );
  dup_2 row_2_d_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:388:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:387:100
    .y     (_row_2_d_x0_1_y),
    .z     (_row_2_d_x0_1_z)
  );
  ADD row_2_n_t1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:389:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_106_2206_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2224:118
    .y     (_row_2_d_x2_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:361:100
    .z     (_row_2_n_t1_1_z)
  );
  MUL row_2_n_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:390:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:353:64
    .y     (_row_2_n_t1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:389:100
    .z     (_row_2_n_x1_1_z)
  );
  dup_2 row_2_d_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:391:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:390:100
    .y     (_row_2_d_x1_1_y),
    .z     (_row_2_d_x1_1_z)
  );
  MUL row_2_n_t2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:392:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_w2_add_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:355:85
    .y     (_row_2_d_x2_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:361:100
    .z     (_row_2_n_t2_1_z)
  );
  SUB row_2_n_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:393:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_d_x1_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:391:100
    .y     (_delay_INT16_71_2204_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2222:114
    .z     (_row_2_n_x2_1_z)
  );
  dup_2 row_2_d_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:394:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:393:100
    .y     (_row_2_d_x2_1_y),
    .z     (_row_2_d_x2_1_z)
  );
  MUL row_2_n_t3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:395:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_w2_sub_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:354:85
    .y     (_delay_INT16_74_2203_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2221:114
    .z     (_row_2_n_t3_1_z)
  );
  ADD row_2_n_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:396:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_d_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:391:100
    .y     (_delay_INT16_188_2202_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2220:118
    .z     (_row_2_n_x3_1_z)
  );
  dup_2 row_2_d_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:397:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:396:100
    .y     (_row_2_d_x3_1_y),
    .z     (_row_2_d_x3_1_z)
  );
  ADD row_2_n_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:398:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_34_2200_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2218:114
    .y     (_row_2_d_x6_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:381:100
    .z     (_row_2_n_x1_2_z)
  );
  dup_2 row_2_d_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:399:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:398:100
    .y     (_row_2_d_x1_2_y),
    .z     (_row_2_d_x1_2_z)
  );
  SUB row_2_n_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:400:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_34_2199_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2217:114
    .y     (_row_2_d_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:381:100
    .z     (_row_2_n_x4_2_z)
  );
  dup_2 row_2_d_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:401:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:400:100
    .y     (_row_2_d_x4_2_y),
    .z     (_row_2_d_x4_2_z)
  );
  ADD row_2_n_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:402:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_143_2198_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2216:118
    .y     (_row_2_d_x7_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:384:100
    .z     (_row_2_n_x6_2_z)
  );
  dup_2 row_2_d_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:403:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:402:100
    .y     (_row_2_d_x6_2_y),
    .z     (_row_2_d_x6_2_z)
  );
  SUB row_2_n_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:404:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_143_2197_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2215:118
    .y     (_row_2_d_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:384:100
    .z     (_row_2_n_x5_2_z)
  );
  dup_2 row_2_d_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:405:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:404:100
    .y     (_row_2_d_x5_2_y),
    .z     (_row_2_d_x5_2_z)
  );
  ADD row_2_n_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:406:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_132_2196_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2214:118
    .y     (_row_2_d_x3_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:397:100
    .z     (_row_2_n_x7_2_z)
  );
  dup_2 row_2_d_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:407:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:406:100
    .y     (_row_2_d_x7_2_y),
    .z     (_row_2_d_x7_2_z)
  );
  SUB row_2_n_x8_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:408:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_132_2317_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2335:118
    .y     (_row_2_d_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:397:100
    .z     (_row_2_n_x8_4_z)
  );
  dup_2 row_2_d_x8_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:409:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x8_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:408:100
    .y     (_row_2_d_x8_4_y),
    .z     (_row_2_d_x8_4_z)
  );
  ADD row_2_n_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:410:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_d_x0_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:388:100
    .y     (_delay_INT16_27_2195_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2213:114
    .z     (_row_2_n_x3_2_z)
  );
  dup_2 row_2_d_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:411:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:410:100
    .y     (_row_2_d_x3_2_y),
    .z     (_row_2_d_x3_2_z)
  );
  SUB row_2_n_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:412:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_d_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:388:100
    .y     (_delay_INT16_27_2192_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2210:114
    .z     (_row_2_n_x0_2_z)
  );
  dup_2 row_2_d_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:413:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:412:100
    .y     (_row_2_d_x0_2_y),
    .z     (_row_2_d_x0_2_z)
  );
  ADD row_2_n_u2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:414:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_72_2191_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2209:114
    .y     (_row_2_d_x5_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:405:100
    .z     (_row_2_n_u2_2_z)
  );
  MUL row_2_n_v2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:415:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_c181_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:345:76
    .y     (_row_2_n_u2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:414:100
    .z     (_row_2_n_v2_2_z)
  );
  ADD row_2_n_w2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:416:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_v2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:415:100
    .y     (_row_2_n_c128_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:343:76
    .z     (_row_2_n_w2_2_z)
  );
  SHR_8 row_2_n_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:417:83
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_w2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:416:100
    .z     (_row_2_n_x2_2_z)
  );
  dup_2 row_2_d_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:418:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:417:83
    .y     (_row_2_d_x2_2_y),
    .z     (_row_2_d_x2_2_z)
  );
  SUB row_2_n_u4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:419:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_72_2188_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2206:114
    .y     (_row_2_d_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:405:100
    .z     (_row_2_n_u4_3_z)
  );
  MUL row_2_n_v4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:420:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_c181_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:346:76
    .y     (_row_2_n_u4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:419:100
    .z     (_row_2_n_v4_3_z)
  );
  ADD row_2_n_w4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:421:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_v4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:420:100
    .y     (_row_2_n_c128_2_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:344:76
    .z     (_row_2_n_w4_3_z)
  );
  SHR_8 row_2_n_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:422:83
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_w4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:421:100
    .z     (_row_2_n_x4_3_z)
  );
  dup_2 row_2_d_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:423:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:422:83
    .y     (_row_2_d_x4_3_y),
    .z     (_row_2_d_x4_3_z)
  );
  ADD row_2_n_tmp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:424:105
    .clock (clock),
    .reset (reset),
    .x     (_row_2_d_x7_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:407:100
    .y     (_delay_INT16_143_2186_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2204:118
    .z     (_row_2_n_tmp_0_z)
  );
  SHR_8 row_2_n_shr_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:425:87
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_tmp_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:424:105
    .z     (_row_2_n_shr_0_z)
  );
  ADD row_2_n_tmp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:426:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_191_2184_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2202:118
    .y     (_row_2_d_x2_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:418:100
    .z     (_row_2_n_tmp_1_z)
  );
  SHR_8 row_2_n_shr_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:427:87
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_tmp_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:426:105
    .z     (_row_2_n_shr_1_z)
  );
  ADD row_2_n_tmp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:428:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_302_2183_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2201:118
    .y     (_row_2_d_x4_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:423:100
    .z     (_row_2_n_tmp_2_z)
  );
  SHR_8 row_2_n_shr_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:429:87
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_tmp_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:428:105
    .z     (_row_2_n_shr_2_z)
  );
  ADD row_2_n_tmp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:430:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_10_2182_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2200:114
    .y     (_row_2_d_x6_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:403:100
    .z     (_row_2_n_tmp_3_z)
  );
  SHR_8 row_2_n_shr_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:431:87
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_tmp_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:430:105
    .z     (_row_2_n_shr_3_z)
  );
  SUB row_2_n_tmp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:432:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_10_2312_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2330:114
    .y     (_row_2_d_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:403:100
    .z     (_row_2_n_tmp_4_z)
  );
  SHR_8 row_2_n_shr_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:433:87
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_tmp_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:432:105
    .z     (_row_2_n_shr_4_z)
  );
  SUB row_2_n_tmp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:434:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_302_2181_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2199:118
    .y     (_row_2_d_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:423:100
    .z     (_row_2_n_tmp_5_z)
  );
  SHR_8 row_2_n_shr_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:435:87
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_tmp_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:434:105
    .z     (_row_2_n_shr_5_z)
  );
  SUB row_2_n_tmp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:436:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_191_2179_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2197:118
    .y     (_row_2_d_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:418:100
    .z     (_row_2_n_tmp_6_z)
  );
  SHR_8 row_2_n_shr_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:437:87
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_tmp_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:436:105
    .z     (_row_2_n_shr_6_z)
  );
  SUB row_2_n_tmp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:438:105
    .clock (clock),
    .reset (reset),
    .x     (_row_2_d_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:407:100
    .y     (_delay_INT16_143_2176_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2194:118
    .z     (_row_2_n_tmp_7_z)
  );
  SHR_8 row_2_n_shr_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:439:87
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_tmp_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:438:105
    .z     (_row_2_n_shr_7_z)
  );
  C128 row_3_n_c128_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:440:76
    .clock (clock),
    .reset (reset),
    .value (_row_3_n_c128_0_value)
  );
  C128 row_3_n_c128_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:441:76
    .clock (clock),
    .reset (reset),
    .value (_row_3_n_c128_1_value)
  );
  C128 row_3_n_c128_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:442:76
    .clock (clock),
    .reset (reset),
    .value (_row_3_n_c128_2_value)
  );
  C181 row_3_n_c181_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:443:76
    .clock (clock),
    .reset (reset),
    .value (_row_3_n_c181_0_value)
  );
  C181 row_3_n_c181_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:444:76
    .clock (clock),
    .reset (reset),
    .value (_row_3_n_c181_1_value)
  );
  W7 row_3_n_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:445:64
    .clock (clock),
    .reset (reset),
    .value (_row_3_n_w7_value)
  );
  W1_sub_W7 row_3_n_w1_sub_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:446:85
    .clock (clock),
    .reset (reset),
    .value (_row_3_n_w1_sub_w7_value)
  );
  W1_add_W7 row_3_n_w1_add_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:447:85
    .clock (clock),
    .reset (reset),
    .value (_row_3_n_w1_add_w7_value)
  );
  W3 row_3_n_w3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:448:64
    .clock (clock),
    .reset (reset),
    .value (_row_3_n_w3_value)
  );
  W3_sub_W5 row_3_n_w3_sub_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:449:85
    .clock (clock),
    .reset (reset),
    .value (_row_3_n_w3_sub_w5_value)
  );
  W3_add_W5 row_3_n_w3_add_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:450:85
    .clock (clock),
    .reset (reset),
    .value (_row_3_n_w3_add_w5_value)
  );
  W6 row_3_n_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:451:64
    .clock (clock),
    .reset (reset),
    .value (_row_3_n_w6_value)
  );
  W2_sub_W6 row_3_n_w2_sub_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:452:85
    .clock (clock),
    .reset (reset),
    .value (_row_3_n_w2_sub_w6_value)
  );
  W2_add_W6 row_3_n_w2_add_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:453:85
    .clock (clock),
    .reset (reset),
    .value (_row_3_n_w2_add_w6_value)
  );
  SHL_11 row_3_n_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:454:83
    .clock (clock),
    .reset (reset),
    .x     (n_in_3_4_x),
    .z     (_row_3_n_x1_0_z)
  );
  SHL_11 row_3_n_t0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:455:83
    .clock (clock),
    .reset (reset),
    .x     (n_in_3_0_x),
    .z     (_row_3_n_t0_0_z)
  );
  ADD row_3_n_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:456:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_t0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:455:83
    .y     (_row_3_n_c128_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:440:76
    .z     (_row_3_n_x0_0_z)
  );
  dup_2 row_3_d_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:457:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:456:100
    .y     (_row_3_d_x0_0_y),
    .z     (_row_3_d_x0_0_z)
  );
  dup_2 row_3_d_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:458:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:454:83
    .y     (_row_3_d_x1_0_y),
    .z     (_row_3_d_x1_0_z)
  );
  dup_2 row_3_d_x2_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:459:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_3_6_x),
    .y     (_row_3_d_x2_0_y),
    .z     (_row_3_d_x2_0_z)
  );
  dup_2 row_3_d_x3_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:460:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_3_2_x),
    .y     (_row_3_d_x3_0_y),
    .z     (_row_3_d_x3_0_z)
  );
  dup_2 row_3_d_x4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:461:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_3_1_x),
    .y     (_row_3_d_x4_0_y),
    .z     (_row_3_d_x4_0_z)
  );
  dup_2 row_3_d_x5_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:462:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_3_7_x),
    .y     (_row_3_d_x5_0_y),
    .z     (_row_3_d_x5_0_z)
  );
  dup_2 row_3_d_x6_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:463:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_3_5_x),
    .y     (_row_3_d_x6_0_y),
    .z     (_row_3_d_x6_0_z)
  );
  dup_2 row_3_d_x7_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:464:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_3_3_x),
    .y     (_row_3_d_x7_0_y),
    .z     (_row_3_d_x7_0_z)
  );
  ADD row_3_n_t8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:465:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_d_x4_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:461:100
    .y     (_delay_INT16_93_2172_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2190:114
    .z     (_row_3_n_t8_1_z)
  );
  MUL row_3_n_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:466:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:445:64
    .y     (_row_3_n_t8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:465:100
    .z     (_row_3_n_x8_1_z)
  );
  dup_2 row_3_d_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:467:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:466:100
    .y     (_row_3_d_x8_1_y),
    .z     (_row_3_d_x8_1_z)
  );
  MUL row_3_n_t4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:468:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_w1_sub_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:446:85
    .y     (_row_3_d_x4_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:461:100
    .z     (_row_3_n_t4_1_z)
  );
  ADD row_3_n_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:469:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_d_x8_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:467:100
    .y     (_delay_INT16_104_2171_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2189:118
    .z     (_row_3_n_x4_1_z)
  );
  dup_2 row_3_d_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:470:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:469:100
    .y     (_row_3_d_x4_1_y),
    .z     (_row_3_d_x4_1_z)
  );
  MUL row_3_n_t5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:471:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_w1_add_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:447:85
    .y     (_delay_INT16_64_2169_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2187:114
    .z     (_row_3_n_t5_1_z)
  );
  SUB row_3_n_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:472:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_d_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:467:100
    .y     (_delay_INT16_53_2168_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2186:114
    .z     (_row_3_n_x5_1_z)
  );
  dup_2 row_3_d_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:473:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:472:100
    .y     (_row_3_d_x5_1_y),
    .z     (_row_3_d_x5_1_z)
  );
  ADD row_3_n_t8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:474:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_d_x6_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:463:100
    .y     (_delay_INT16_60_2167_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2185:114
    .z     (_row_3_n_t8_2_z)
  );
  MUL row_3_n_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:475:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_w3_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:448:64
    .y     (_row_3_n_t8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:474:100
    .z     (_row_3_n_x8_2_z)
  );
  dup_2 row_3_d_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:476:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:475:100
    .y     (_row_3_d_x8_2_y),
    .z     (_row_3_d_x8_2_z)
  );
  MUL row_3_n_t6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:477:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_w3_sub_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:449:85
    .y     (_row_3_d_x6_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:463:100
    .z     (_row_3_n_t6_1_z)
  );
  SUB row_3_n_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:478:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_d_x8_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:476:100
    .y     (_delay_INT16_74_2175_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2193:114
    .z     (_row_3_n_x6_1_z)
  );
  dup_2 row_3_d_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:479:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:478:100
    .y     (_row_3_d_x6_1_y),
    .z     (_row_3_d_x6_1_z)
  );
  MUL row_3_n_t7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:480:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_w3_add_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:450:85
    .y     (_delay_INT16_11_2166_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2184:114
    .z     (_row_3_n_t7_1_z)
  );
  SUB row_3_n_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:481:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_d_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:476:100
    .y     (_delay_INT16_206_2164_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2182:118
    .z     (_row_3_n_x7_1_z)
  );
  dup_2 row_3_d_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:482:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:481:100
    .y     (_row_3_d_x7_1_y),
    .z     (_row_3_d_x7_1_z)
  );
  ADD row_3_n_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:483:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_d_x0_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:457:100
    .y     (_delay_INT16_180_2194_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2212:118
    .z     (_row_3_n_x8_3_z)
  );
  dup_2 row_3_d_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:484:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:483:100
    .y     (_row_3_d_x8_3_y),
    .z     (_row_3_d_x8_3_z)
  );
  SUB row_3_n_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:485:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_d_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:457:100
    .y     (_delay_INT16_180_2218_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2236:118
    .z     (_row_3_n_x0_1_z)
  );
  dup_2 row_3_d_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:486:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:485:100
    .y     (_row_3_d_x0_1_y),
    .z     (_row_3_d_x0_1_z)
  );
  ADD row_3_n_t1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:487:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_d_x3_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:460:100
    .y     (_delay_INT16_96_2163_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2181:114
    .z     (_row_3_n_t1_1_z)
  );
  MUL row_3_n_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:488:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:451:64
    .y     (_row_3_n_t1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:487:100
    .z     (_row_3_n_x1_1_z)
  );
  dup_2 row_3_d_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:489:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:488:100
    .y     (_row_3_d_x1_1_y),
    .z     (_row_3_d_x1_1_z)
  );
  MUL row_3_n_t2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:490:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_w2_add_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:453:85
    .y     (_row_3_d_x2_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:459:100
    .z     (_row_3_n_t2_1_z)
  );
  SUB row_3_n_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:491:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_d_x1_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:489:100
    .y     (_delay_INT16_289_2212_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2230:118
    .z     (_row_3_n_x2_1_z)
  );
  dup_2 row_3_d_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:492:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:491:100
    .y     (_row_3_d_x2_1_y),
    .z     (_row_3_d_x2_1_z)
  );
  MUL row_3_n_t3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:493:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_w2_sub_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:452:85
    .y     (_row_3_d_x3_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:460:100
    .z     (_row_3_n_t3_1_z)
  );
  ADD row_3_n_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:494:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_d_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:489:100
    .y     (_delay_INT16_108_2298_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2316:118
    .z     (_row_3_n_x3_1_z)
  );
  dup_2 row_3_d_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:495:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:494:100
    .y     (_row_3_d_x3_1_y),
    .z     (_row_3_d_x3_1_z)
  );
  ADD row_3_n_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:496:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_11_2162_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2180:114
    .y     (_row_3_d_x6_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:479:100
    .z     (_row_3_n_x1_2_z)
  );
  dup_2 row_3_d_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:497:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:496:100
    .y     (_row_3_d_x1_2_y),
    .z     (_row_3_d_x1_2_z)
  );
  SUB row_3_n_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:498:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_11_2161_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2179:114
    .y     (_row_3_d_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:479:100
    .z     (_row_3_n_x4_2_z)
  );
  dup_2 row_3_d_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:499:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:498:100
    .y     (_row_3_d_x4_2_y),
    .z     (_row_3_d_x4_2_z)
  );
  ADD row_3_n_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:500:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_49_2160_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2178:114
    .y     (_row_3_d_x7_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:482:100
    .z     (_row_3_n_x6_2_z)
  );
  dup_2 row_3_d_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:501:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:500:100
    .y     (_row_3_d_x6_2_y),
    .z     (_row_3_d_x6_2_z)
  );
  SUB row_3_n_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:502:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_49_2159_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2177:114
    .y     (_row_3_d_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:482:100
    .z     (_row_3_n_x5_2_z)
  );
  dup_2 row_3_d_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:503:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:502:100
    .y     (_row_3_d_x5_2_y),
    .z     (_row_3_d_x5_2_z)
  );
  ADD row_3_n_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:504:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_109_2223_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2241:118
    .y     (_row_3_d_x3_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:495:100
    .z     (_row_3_n_x7_2_z)
  );
  dup_2 row_3_d_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:505:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:504:100
    .y     (_row_3_d_x7_2_y),
    .z     (_row_3_d_x7_2_z)
  );
  SUB row_3_n_x8_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:506:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_109_2207_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2225:118
    .y     (_row_3_d_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:495:100
    .z     (_row_3_n_x8_4_z)
  );
  dup_2 row_3_d_x8_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:507:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x8_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:506:100
    .y     (_row_3_d_x8_4_y),
    .z     (_row_3_d_x8_4_z)
  );
  ADD row_3_n_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:508:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_40_2170_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2188:114
    .y     (_row_3_d_x2_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:492:100
    .z     (_row_3_n_x3_2_z)
  );
  dup_2 row_3_d_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:509:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:508:100
    .y     (_row_3_d_x3_2_y),
    .z     (_row_3_d_x3_2_z)
  );
  SUB row_3_n_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:510:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_40_2157_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2175:114
    .y     (_row_3_d_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:492:100
    .z     (_row_3_n_x0_2_z)
  );
  dup_2 row_3_d_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:511:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:510:100
    .y     (_row_3_d_x0_2_y),
    .z     (_row_3_d_x0_2_z)
  );
  ADD row_3_n_u2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:512:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_125_2155_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2173:118
    .y     (_row_3_d_x5_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:503:100
    .z     (_row_3_n_u2_2_z)
  );
  MUL row_3_n_v2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:513:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_c181_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:443:76
    .y     (_row_3_n_u2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:512:100
    .z     (_row_3_n_v2_2_z)
  );
  ADD row_3_n_w2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:514:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_v2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:513:100
    .y     (_row_3_n_c128_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:441:76
    .z     (_row_3_n_w2_2_z)
  );
  SHR_8 row_3_n_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:515:83
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_w2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:514:100
    .z     (_row_3_n_x2_2_z)
  );
  dup_2 row_3_d_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:516:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:515:83
    .y     (_row_3_d_x2_2_y),
    .z     (_row_3_d_x2_2_z)
  );
  SUB row_3_n_u4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:517:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_125_2154_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2172:118
    .y     (_row_3_d_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:503:100
    .z     (_row_3_n_u4_3_z)
  );
  MUL row_3_n_v4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:518:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_c181_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:444:76
    .y     (_row_3_n_u4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:517:100
    .z     (_row_3_n_v4_3_z)
  );
  ADD row_3_n_w4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:519:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_v4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:518:100
    .y     (_row_3_n_c128_2_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:442:76
    .z     (_row_3_n_w4_3_z)
  );
  SHR_8 row_3_n_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:520:83
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_w4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:519:100
    .z     (_row_3_n_x4_3_z)
  );
  dup_2 row_3_d_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:521:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:520:83
    .y     (_row_3_d_x4_3_y),
    .z     (_row_3_d_x4_3_z)
  );
  ADD row_3_n_tmp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:522:105
    .clock (clock),
    .reset (reset),
    .x     (_row_3_d_x7_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:505:100
    .y     (_delay_INT16_127_2153_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2171:118
    .z     (_row_3_n_tmp_0_z)
  );
  SHR_8 row_3_n_shr_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:523:87
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_tmp_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:522:105
    .z     (_row_3_n_shr_0_z)
  );
  ADD row_3_n_tmp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:524:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_157_2152_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2170:118
    .y     (_row_3_d_x2_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:516:100
    .z     (_row_3_n_tmp_1_z)
  );
  SHR_8 row_3_n_shr_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:525:87
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_tmp_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:524:105
    .z     (_row_3_n_shr_1_z)
  );
  ADD row_3_n_tmp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:526:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_152_2307_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2325:118
    .y     (_row_3_d_x4_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:521:100
    .z     (_row_3_n_tmp_2_z)
  );
  SHR_8 row_3_n_shr_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:527:87
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_tmp_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:526:105
    .z     (_row_3_n_shr_2_z)
  );
  ADD row_3_n_tmp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:528:105
    .clock (clock),
    .reset (reset),
    .x     (_row_3_d_x8_4_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:507:100
    .y     (_delay_INT16_31_2150_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2168:114
    .z     (_row_3_n_tmp_3_z)
  );
  SHR_8 row_3_n_shr_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:529:87
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_tmp_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:528:105
    .z     (_row_3_n_shr_3_z)
  );
  SUB row_3_n_tmp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:530:105
    .clock (clock),
    .reset (reset),
    .x     (_row_3_d_x8_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:507:100
    .y     (_delay_INT16_31_2280_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2298:114
    .z     (_row_3_n_tmp_4_z)
  );
  SHR_8 row_3_n_shr_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:531:87
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_tmp_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:530:105
    .z     (_row_3_n_shr_4_z)
  );
  SUB row_3_n_tmp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:532:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_152_2149_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2167:118
    .y     (_row_3_d_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:521:100
    .z     (_row_3_n_tmp_5_z)
  );
  SHR_8 row_3_n_shr_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:533:87
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_tmp_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:532:105
    .z     (_row_3_n_shr_5_z)
  );
  SUB row_3_n_tmp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:534:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_157_2148_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2166:118
    .y     (_row_3_d_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:516:100
    .z     (_row_3_n_tmp_6_z)
  );
  SHR_8 row_3_n_shr_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:535:87
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_tmp_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:534:105
    .z     (_row_3_n_shr_6_z)
  );
  SUB row_3_n_tmp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:536:105
    .clock (clock),
    .reset (reset),
    .x     (_row_3_d_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:505:100
    .y     (_delay_INT16_127_2147_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2165:118
    .z     (_row_3_n_tmp_7_z)
  );
  SHR_8 row_3_n_shr_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:537:87
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_tmp_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:536:105
    .z     (_row_3_n_shr_7_z)
  );
  C128 row_4_n_c128_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:538:76
    .clock (clock),
    .reset (reset),
    .value (_row_4_n_c128_0_value)
  );
  C128 row_4_n_c128_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:539:76
    .clock (clock),
    .reset (reset),
    .value (_row_4_n_c128_1_value)
  );
  C128 row_4_n_c128_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:540:76
    .clock (clock),
    .reset (reset),
    .value (_row_4_n_c128_2_value)
  );
  C181 row_4_n_c181_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:541:76
    .clock (clock),
    .reset (reset),
    .value (_row_4_n_c181_0_value)
  );
  C181 row_4_n_c181_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:542:76
    .clock (clock),
    .reset (reset),
    .value (_row_4_n_c181_1_value)
  );
  W7 row_4_n_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:543:64
    .clock (clock),
    .reset (reset),
    .value (_row_4_n_w7_value)
  );
  W1_sub_W7 row_4_n_w1_sub_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:544:85
    .clock (clock),
    .reset (reset),
    .value (_row_4_n_w1_sub_w7_value)
  );
  W1_add_W7 row_4_n_w1_add_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:545:85
    .clock (clock),
    .reset (reset),
    .value (_row_4_n_w1_add_w7_value)
  );
  W3 row_4_n_w3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:546:64
    .clock (clock),
    .reset (reset),
    .value (_row_4_n_w3_value)
  );
  W3_sub_W5 row_4_n_w3_sub_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:547:85
    .clock (clock),
    .reset (reset),
    .value (_row_4_n_w3_sub_w5_value)
  );
  W3_add_W5 row_4_n_w3_add_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:548:85
    .clock (clock),
    .reset (reset),
    .value (_row_4_n_w3_add_w5_value)
  );
  W6 row_4_n_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:549:64
    .clock (clock),
    .reset (reset),
    .value (_row_4_n_w6_value)
  );
  W2_sub_W6 row_4_n_w2_sub_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:550:85
    .clock (clock),
    .reset (reset),
    .value (_row_4_n_w2_sub_w6_value)
  );
  W2_add_W6 row_4_n_w2_add_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:551:85
    .clock (clock),
    .reset (reset),
    .value (_row_4_n_w2_add_w6_value)
  );
  SHL_11 row_4_n_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:552:83
    .clock (clock),
    .reset (reset),
    .x     (n_in_4_4_x),
    .z     (_row_4_n_x1_0_z)
  );
  SHL_11 row_4_n_t0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:553:83
    .clock (clock),
    .reset (reset),
    .x     (n_in_4_0_x),
    .z     (_row_4_n_t0_0_z)
  );
  ADD row_4_n_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:554:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_t0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:553:83
    .y     (_row_4_n_c128_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:538:76
    .z     (_row_4_n_x0_0_z)
  );
  dup_2 row_4_d_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:555:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:554:100
    .y     (_row_4_d_x0_0_y),
    .z     (_row_4_d_x0_0_z)
  );
  dup_2 row_4_d_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:556:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:552:83
    .y     (_row_4_d_x1_0_y),
    .z     (_row_4_d_x1_0_z)
  );
  dup_2 row_4_d_x2_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:557:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_4_6_x),
    .y     (_row_4_d_x2_0_y),
    .z     (_row_4_d_x2_0_z)
  );
  dup_2 row_4_d_x3_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:558:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_4_2_x),
    .y     (_row_4_d_x3_0_y),
    .z     (_row_4_d_x3_0_z)
  );
  dup_2 row_4_d_x4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:559:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_4_1_x),
    .y     (_row_4_d_x4_0_y),
    .z     (_row_4_d_x4_0_z)
  );
  dup_2 row_4_d_x5_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:560:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_4_7_x),
    .y     (_row_4_d_x5_0_y),
    .z     (_row_4_d_x5_0_z)
  );
  dup_2 row_4_d_x6_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:561:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_4_5_x),
    .y     (_row_4_d_x6_0_y),
    .z     (_row_4_d_x6_0_z)
  );
  dup_2 row_4_d_x7_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:562:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_4_3_x),
    .y     (_row_4_d_x7_0_y),
    .z     (_row_4_d_x7_0_z)
  );
  ADD row_4_n_t8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:563:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_60_2143_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2161:114
    .y     (_row_4_d_x5_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:560:100
    .z     (_row_4_n_t8_1_z)
  );
  MUL row_4_n_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:564:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:543:64
    .y     (_row_4_n_t8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:563:100
    .z     (_row_4_n_x8_1_z)
  );
  dup_2 row_4_d_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:565:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:564:100
    .y     (_row_4_d_x8_1_y),
    .z     (_row_4_d_x8_1_z)
  );
  MUL row_4_n_t4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:566:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_w1_sub_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:544:85
    .y     (_delay_INT16_28_2141_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2159:114
    .z     (_row_4_n_t4_1_z)
  );
  ADD row_4_n_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:567:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_d_x8_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:565:100
    .y     (_delay_INT16_268_2299_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2317:118
    .z     (_row_4_n_x4_1_z)
  );
  dup_2 row_4_d_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:568:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:567:100
    .y     (_row_4_d_x4_1_y),
    .z     (_row_4_d_x4_1_z)
  );
  MUL row_4_n_t5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:569:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_w1_add_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:545:85
    .y     (_row_4_d_x5_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:560:100
    .z     (_row_4_n_t5_1_z)
  );
  SUB row_4_n_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:570:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_d_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:565:100
    .y     (_delay_INT16_230_2308_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2326:118
    .z     (_row_4_n_x5_1_z)
  );
  dup_2 row_4_d_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:571:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:570:100
    .y     (_row_4_d_x5_1_y),
    .z     (_row_4_d_x5_1_z)
  );
  ADD row_4_n_t8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:572:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_d_x6_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:561:100
    .y     (_delay_INT16_24_2140_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2158:114
    .z     (_row_4_n_t8_2_z)
  );
  MUL row_4_n_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:573:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_w3_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:546:64
    .y     (_row_4_n_t8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:572:100
    .z     (_row_4_n_x8_2_z)
  );
  dup_2 row_4_d_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:574:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:573:100
    .y     (_row_4_d_x8_2_y),
    .z     (_row_4_d_x8_2_z)
  );
  MUL row_4_n_t6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:575:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_w3_sub_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:547:85
    .y     (_row_4_d_x6_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:561:100
    .z     (_row_4_n_t6_1_z)
  );
  SUB row_4_n_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:576:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_d_x8_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:574:100
    .y     (_delay_INT16_131_2139_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2157:118
    .z     (_row_4_n_x6_1_z)
  );
  dup_2 row_4_d_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:577:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:576:100
    .y     (_row_4_d_x6_1_y),
    .z     (_row_4_d_x6_1_z)
  );
  MUL row_4_n_t7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:578:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_w3_add_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:548:85
    .y     (_row_4_d_x7_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:562:100
    .z     (_row_4_n_t7_1_z)
  );
  SUB row_4_n_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:579:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_d_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:574:100
    .y     (_delay_INT16_234_2318_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2336:118
    .z     (_row_4_n_x7_1_z)
  );
  dup_2 row_4_d_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:580:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:579:100
    .y     (_row_4_d_x7_1_y),
    .z     (_row_4_d_x7_1_z)
  );
  ADD row_4_n_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:581:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_d_x0_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:555:100
    .y     (_delay_INT16_184_2136_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2154:118
    .z     (_row_4_n_x8_3_z)
  );
  dup_2 row_4_d_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:582:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:581:100
    .y     (_row_4_d_x8_3_y),
    .z     (_row_4_d_x8_3_z)
  );
  SUB row_4_n_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:583:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_d_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:555:100
    .y     (_delay_INT16_184_2187_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2205:118
    .z     (_row_4_n_x0_1_z)
  );
  dup_2 row_4_d_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:584:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:583:100
    .y     (_row_4_d_x0_1_y),
    .z     (_row_4_d_x0_1_z)
  );
  ADD row_4_n_t1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:585:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_72_2259_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2277:114
    .y     (_row_4_d_x2_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:557:100
    .z     (_row_4_n_t1_1_z)
  );
  MUL row_4_n_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:586:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:549:64
    .y     (_row_4_n_t1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:585:100
    .z     (_row_4_n_x1_1_z)
  );
  dup_2 row_4_d_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:587:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:586:100
    .y     (_row_4_d_x1_1_y),
    .z     (_row_4_d_x1_1_z)
  );
  MUL row_4_n_t2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:588:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_w2_add_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:551:85
    .y     (_row_4_d_x2_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:557:100
    .z     (_row_4_n_t2_1_z)
  );
  SUB row_4_n_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:589:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_d_x1_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:587:100
    .y     (_delay_INT16_145_2134_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2152:118
    .z     (_row_4_n_x2_1_z)
  );
  dup_2 row_4_d_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:590:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:589:100
    .y     (_row_4_d_x2_1_y),
    .z     (_row_4_d_x2_1_z)
  );
  MUL row_4_n_t3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:591:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_w2_sub_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:550:85
    .y     (_row_4_d_x3_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:558:100
    .z     (_row_4_n_t3_1_z)
  );
  ADD row_4_n_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:592:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_d_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:587:100
    .y     (_delay_INT16_248_2145_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2163:118
    .z     (_row_4_n_x3_1_z)
  );
  dup_2 row_4_d_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:593:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:592:100
    .y     (_row_4_d_x3_1_y),
    .z     (_row_4_d_x3_1_z)
  );
  ADD row_4_n_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:594:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_79_2132_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2150:114
    .y     (_row_4_d_x6_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:577:100
    .z     (_row_4_n_x1_2_z)
  );
  dup_2 row_4_d_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:595:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:594:100
    .y     (_row_4_d_x1_2_y),
    .z     (_row_4_d_x1_2_z)
  );
  SUB row_4_n_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:596:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_79_2131_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2149:114
    .y     (_row_4_d_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:577:100
    .z     (_row_4_n_x4_2_z)
  );
  dup_2 row_4_d_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:597:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:596:100
    .y     (_row_4_d_x4_2_y),
    .z     (_row_4_d_x4_2_z)
  );
  ADD row_4_n_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:598:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_95_2130_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2148:114
    .y     (_row_4_d_x7_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:580:100
    .z     (_row_4_n_x6_2_z)
  );
  dup_2 row_4_d_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:599:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:598:100
    .y     (_row_4_d_x6_2_y),
    .z     (_row_4_d_x6_2_z)
  );
  SUB row_4_n_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:600:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_95_2129_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2147:114
    .y     (_row_4_d_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:580:100
    .z     (_row_4_n_x5_2_z)
  );
  dup_2 row_4_d_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:601:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:600:100
    .y     (_row_4_d_x5_2_y),
    .z     (_row_4_d_x5_2_z)
  );
  ADD row_4_n_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:602:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_229_2128_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2146:118
    .y     (_row_4_d_x3_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:593:100
    .z     (_row_4_n_x7_2_z)
  );
  dup_2 row_4_d_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:603:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:602:100
    .y     (_row_4_d_x7_2_y),
    .z     (_row_4_d_x7_2_z)
  );
  SUB row_4_n_x8_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:604:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_229_2126_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2144:118
    .y     (_row_4_d_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:593:100
    .z     (_row_4_n_x8_4_z)
  );
  dup_2 row_4_d_x8_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:605:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x8_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:604:100
    .y     (_row_4_d_x8_4_y),
    .z     (_row_4_d_x8_4_z)
  );
  ADD row_4_n_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:606:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_166_2125_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2143:118
    .y     (_row_4_d_x2_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:590:100
    .z     (_row_4_n_x3_2_z)
  );
  dup_2 row_4_d_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:607:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:606:100
    .y     (_row_4_d_x3_2_y),
    .z     (_row_4_d_x3_2_z)
  );
  SUB row_4_n_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:608:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_166_2124_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2142:118
    .y     (_row_4_d_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:590:100
    .z     (_row_4_n_x0_2_z)
  );
  dup_2 row_4_d_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:609:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:608:100
    .y     (_row_4_d_x0_2_y),
    .z     (_row_4_d_x0_2_z)
  );
  ADD row_4_n_u2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:610:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_114_2122_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2140:118
    .y     (_row_4_d_x5_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:601:100
    .z     (_row_4_n_u2_2_z)
  );
  MUL row_4_n_v2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:611:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_c181_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:541:76
    .y     (_row_4_n_u2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:610:100
    .z     (_row_4_n_v2_2_z)
  );
  ADD row_4_n_w2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:612:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_v2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:611:100
    .y     (_row_4_n_c128_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:539:76
    .z     (_row_4_n_w2_2_z)
  );
  SHR_8 row_4_n_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:613:83
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_w2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:612:100
    .z     (_row_4_n_x2_2_z)
  );
  dup_2 row_4_d_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:614:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:613:83
    .y     (_row_4_d_x2_2_y),
    .z     (_row_4_d_x2_2_z)
  );
  SUB row_4_n_u4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:615:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_114_2120_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2138:118
    .y     (_row_4_d_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:601:100
    .z     (_row_4_n_u4_3_z)
  );
  MUL row_4_n_v4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:616:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_c181_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:542:76
    .y     (_row_4_n_u4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:615:100
    .z     (_row_4_n_v4_3_z)
  );
  ADD row_4_n_w4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:617:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_v4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:616:100
    .y     (_row_4_n_c128_2_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:540:76
    .z     (_row_4_n_w4_3_z)
  );
  SHR_8 row_4_n_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:618:83
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_w4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:617:100
    .z     (_row_4_n_x4_3_z)
  );
  dup_2 row_4_d_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:619:100
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:618:83
    .y     (_row_4_d_x4_3_y),
    .z     (_row_4_d_x4_3_z)
  );
  ADD row_4_n_tmp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:620:105
    .clock (clock),
    .reset (reset),
    .x     (_row_4_d_x7_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:603:100
    .y     (_delay_INT16_83_2119_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2137:114
    .z     (_row_4_n_tmp_0_z)
  );
  SHR_8 row_4_n_shr_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:621:87
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_tmp_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:620:105
    .z     (_row_4_n_shr_0_z)
  );
  ADD row_4_n_tmp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:622:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_248_2118_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2136:118
    .y     (_row_4_d_x2_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:614:100
    .z     (_row_4_n_tmp_1_z)
  );
  SHR_8 row_4_n_shr_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:623:87
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_tmp_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:622:105
    .z     (_row_4_n_shr_1_z)
  );
  ADD row_4_n_tmp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:624:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_350_2117_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2135:118
    .y     (_row_4_d_x4_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:619:100
    .z     (_row_4_n_tmp_2_z)
  );
  SHR_8 row_4_n_shr_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:625:87
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_tmp_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:624:105
    .z     (_row_4_n_shr_2_z)
  );
  ADD row_4_n_tmp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:626:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_58_2325_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2343:114
    .y     (_row_4_d_x6_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:599:100
    .z     (_row_4_n_tmp_3_z)
  );
  SHR_8 row_4_n_shr_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:627:87
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_tmp_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:626:105
    .z     (_row_4_n_shr_3_z)
  );
  SUB row_4_n_tmp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:628:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_58_2217_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2235:114
    .y     (_row_4_d_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:599:100
    .z     (_row_4_n_tmp_4_z)
  );
  SHR_8 row_4_n_shr_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:629:87
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_tmp_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:628:105
    .z     (_row_4_n_shr_4_z)
  );
  SUB row_4_n_tmp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:630:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_350_2284_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2302:118
    .y     (_row_4_d_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:619:100
    .z     (_row_4_n_tmp_5_z)
  );
  SHR_8 row_4_n_shr_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:631:87
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_tmp_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:630:105
    .z     (_row_4_n_shr_5_z)
  );
  SUB row_4_n_tmp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:632:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_248_2114_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2132:118
    .y     (_row_4_d_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:614:100
    .z     (_row_4_n_tmp_6_z)
  );
  SHR_8 row_4_n_shr_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:633:87
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_tmp_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:632:105
    .z     (_row_4_n_shr_6_z)
  );
  SUB row_4_n_tmp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:634:105
    .clock (clock),
    .reset (reset),
    .x     (_row_4_d_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:603:100
    .y     (_delay_INT16_83_2113_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2131:114
    .z     (_row_4_n_tmp_7_z)
  );
  SHR_8 row_4_n_shr_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:635:87
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_tmp_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:634:105
    .z     (_row_4_n_shr_7_z)
  );
  C128 row_5_n_c128_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:636:76
    .clock (clock),
    .reset (reset),
    .value (_row_5_n_c128_0_value)
  );
  C128 row_5_n_c128_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:637:76
    .clock (clock),
    .reset (reset),
    .value (_row_5_n_c128_1_value)
  );
  C128 row_5_n_c128_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:638:76
    .clock (clock),
    .reset (reset),
    .value (_row_5_n_c128_2_value)
  );
  C181 row_5_n_c181_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:639:76
    .clock (clock),
    .reset (reset),
    .value (_row_5_n_c181_0_value)
  );
  C181 row_5_n_c181_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:640:76
    .clock (clock),
    .reset (reset),
    .value (_row_5_n_c181_1_value)
  );
  W7 row_5_n_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:641:64
    .clock (clock),
    .reset (reset),
    .value (_row_5_n_w7_value)
  );
  W1_sub_W7 row_5_n_w1_sub_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:642:85
    .clock (clock),
    .reset (reset),
    .value (_row_5_n_w1_sub_w7_value)
  );
  W1_add_W7 row_5_n_w1_add_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:643:85
    .clock (clock),
    .reset (reset),
    .value (_row_5_n_w1_add_w7_value)
  );
  W3 row_5_n_w3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:644:64
    .clock (clock),
    .reset (reset),
    .value (_row_5_n_w3_value)
  );
  W3_sub_W5 row_5_n_w3_sub_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:645:85
    .clock (clock),
    .reset (reset),
    .value (_row_5_n_w3_sub_w5_value)
  );
  W3_add_W5 row_5_n_w3_add_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:646:85
    .clock (clock),
    .reset (reset),
    .value (_row_5_n_w3_add_w5_value)
  );
  W6 row_5_n_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:647:64
    .clock (clock),
    .reset (reset),
    .value (_row_5_n_w6_value)
  );
  W2_sub_W6 row_5_n_w2_sub_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:648:85
    .clock (clock),
    .reset (reset),
    .value (_row_5_n_w2_sub_w6_value)
  );
  W2_add_W6 row_5_n_w2_add_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:649:85
    .clock (clock),
    .reset (reset),
    .value (_row_5_n_w2_add_w6_value)
  );
  SHL_11 row_5_n_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:650:83
    .clock (clock),
    .reset (reset),
    .x     (n_in_5_4_x),
    .z     (_row_5_n_x1_0_z)
  );
  SHL_11 row_5_n_t0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:651:83
    .clock (clock),
    .reset (reset),
    .x     (n_in_5_0_x),
    .z     (_row_5_n_t0_0_z)
  );
  ADD row_5_n_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:652:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_t0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:651:83
    .y     (_row_5_n_c128_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:636:76
    .z     (_row_5_n_x0_0_z)
  );
  dup_2 row_5_d_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:653:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:652:100
    .y     (_row_5_d_x0_0_y),
    .z     (_row_5_d_x0_0_z)
  );
  dup_2 row_5_d_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:654:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:650:83
    .y     (_row_5_d_x1_0_y),
    .z     (_row_5_d_x1_0_z)
  );
  dup_2 row_5_d_x2_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:655:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_5_6_x),
    .y     (_row_5_d_x2_0_y),
    .z     (_row_5_d_x2_0_z)
  );
  dup_2 row_5_d_x3_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:656:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_5_2_x),
    .y     (_row_5_d_x3_0_y),
    .z     (_row_5_d_x3_0_z)
  );
  dup_2 row_5_d_x4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:657:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_5_1_x),
    .y     (_row_5_d_x4_0_y),
    .z     (_row_5_d_x4_0_z)
  );
  dup_2 row_5_d_x5_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:658:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_5_7_x),
    .y     (_row_5_d_x5_0_y),
    .z     (_row_5_d_x5_0_z)
  );
  dup_2 row_5_d_x6_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:659:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_5_5_x),
    .y     (_row_5_d_x6_0_y),
    .z     (_row_5_d_x6_0_z)
  );
  dup_2 row_5_d_x7_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:660:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_5_3_x),
    .y     (_row_5_d_x7_0_y),
    .z     (_row_5_d_x7_0_z)
  );
  ADD row_5_n_t8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:661:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_d_x4_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:657:100
    .y     (_delay_INT16_87_2110_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2128:114
    .z     (_row_5_n_t8_1_z)
  );
  MUL row_5_n_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:662:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:641:64
    .y     (_row_5_n_t8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:661:100
    .z     (_row_5_n_x8_1_z)
  );
  dup_2 row_5_d_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:663:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:662:100
    .y     (_row_5_d_x8_1_y),
    .z     (_row_5_d_x8_1_z)
  );
  MUL row_5_n_t4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:664:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_w1_sub_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:642:85
    .y     (_row_5_d_x4_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:657:100
    .z     (_row_5_n_t4_1_z)
  );
  ADD row_5_n_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:665:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_d_x8_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:663:100
    .y     (_delay_INT16_10_2109_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2127:114
    .z     (_row_5_n_x4_1_z)
  );
  dup_2 row_5_d_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:666:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:665:100
    .y     (_row_5_d_x4_1_y),
    .z     (_row_5_d_x4_1_z)
  );
  MUL row_5_n_t5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:667:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_w1_add_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:643:85
    .y     (_delay_INT16_13_2108_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2126:114
    .z     (_row_5_n_t5_1_z)
  );
  SUB row_5_n_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:668:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_d_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:663:100
    .y     (_delay_INT16_121_2107_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2125:118
    .z     (_row_5_n_x5_1_z)
  );
  dup_2 row_5_d_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:669:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:668:100
    .y     (_row_5_d_x5_1_y),
    .z     (_row_5_d_x5_1_z)
  );
  ADD row_5_n_t8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:670:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_d_x6_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:659:100
    .y     (_delay_INT16_10_2106_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2124:114
    .z     (_row_5_n_t8_2_z)
  );
  MUL row_5_n_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:671:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_w3_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:644:64
    .y     (_row_5_n_t8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:670:100
    .z     (_row_5_n_x8_2_z)
  );
  dup_2 row_5_d_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:672:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:671:100
    .y     (_row_5_d_x8_2_y),
    .z     (_row_5_d_x8_2_z)
  );
  MUL row_5_n_t6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:673:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_w3_sub_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:645:85
    .y     (_row_5_d_x6_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:659:100
    .z     (_row_5_n_t6_1_z)
  );
  SUB row_5_n_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:674:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_d_x8_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:672:100
    .y     (_delay_INT16_43_2105_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2123:114
    .z     (_row_5_n_x6_1_z)
  );
  dup_2 row_5_d_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:675:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:674:100
    .y     (_row_5_d_x6_1_y),
    .z     (_row_5_d_x6_1_z)
  );
  MUL row_5_n_t7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:676:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_w3_add_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:646:85
    .y     (_row_5_d_x7_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:660:100
    .z     (_row_5_n_t7_1_z)
  );
  SUB row_5_n_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:677:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_d_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:672:100
    .y     (_delay_INT16_87_2104_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2122:114
    .z     (_row_5_n_x7_1_z)
  );
  dup_2 row_5_d_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:678:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:677:100
    .y     (_row_5_d_x7_1_y),
    .z     (_row_5_d_x7_1_z)
  );
  ADD row_5_n_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:679:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_8_2103_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2121:110
    .y     (_row_5_d_x1_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:654:100
    .z     (_row_5_n_x8_3_z)
  );
  dup_2 row_5_d_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:680:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:679:100
    .y     (_row_5_d_x8_3_y),
    .z     (_row_5_d_x8_3_z)
  );
  SUB row_5_n_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:681:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_8_2102_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2120:110
    .y     (_row_5_d_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:654:100
    .z     (_row_5_n_x0_1_z)
  );
  dup_2 row_5_d_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:682:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:681:100
    .y     (_row_5_d_x0_1_y),
    .z     (_row_5_d_x0_1_z)
  );
  ADD row_5_n_t1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:683:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_d_x3_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:656:100
    .y     (_delay_INT16_31_2101_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2119:114
    .z     (_row_5_n_t1_1_z)
  );
  MUL row_5_n_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:684:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:647:64
    .y     (_row_5_n_t1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:683:100
    .z     (_row_5_n_x1_1_z)
  );
  dup_2 row_5_d_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:685:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:684:100
    .y     (_row_5_d_x1_1_y),
    .z     (_row_5_d_x1_1_z)
  );
  MUL row_5_n_t2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:686:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_w2_add_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:649:85
    .y     (_row_5_d_x2_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:655:100
    .z     (_row_5_n_t2_1_z)
  );
  SUB row_5_n_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:687:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_d_x1_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:685:100
    .y     (_delay_INT16_226_2100_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2118:118
    .z     (_row_5_n_x2_1_z)
  );
  dup_2 row_5_d_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:688:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:687:100
    .y     (_row_5_d_x2_1_y),
    .z     (_row_5_d_x2_1_z)
  );
  MUL row_5_n_t3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:689:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_w2_sub_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:648:85
    .y     (_row_5_d_x3_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:656:100
    .z     (_row_5_n_t3_1_z)
  );
  ADD row_5_n_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:690:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_d_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:685:100
    .y     (_delay_INT16_224_2099_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2117:118
    .z     (_row_5_n_x3_1_z)
  );
  dup_2 row_5_d_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:691:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:690:100
    .y     (_row_5_d_x3_1_y),
    .z     (_row_5_d_x3_1_z)
  );
  ADD row_5_n_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:692:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_d_x4_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:666:100
    .y     (_delay_INT16_5_2098_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2116:110
    .z     (_row_5_n_x1_2_z)
  );
  dup_2 row_5_d_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:693:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:692:100
    .y     (_row_5_d_x1_2_y),
    .z     (_row_5_d_x1_2_z)
  );
  SUB row_5_n_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:694:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_d_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:666:100
    .y     (_delay_INT16_5_2096_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2114:110
    .z     (_row_5_n_x4_2_z)
  );
  dup_2 row_5_d_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:695:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:694:100
    .y     (_row_5_d_x4_2_y),
    .z     (_row_5_d_x4_2_z)
  );
  ADD row_5_n_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:696:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_d_x5_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:669:100
    .y     (_delay_INT16_61_2095_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2113:114
    .z     (_row_5_n_x6_2_z)
  );
  dup_2 row_5_d_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:697:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:696:100
    .y     (_row_5_d_x6_2_y),
    .z     (_row_5_d_x6_2_z)
  );
  SUB row_5_n_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:698:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_d_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:669:100
    .y     (_delay_INT16_61_2094_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2112:114
    .z     (_row_5_n_x5_2_z)
  );
  dup_2 row_5_d_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:699:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:698:100
    .y     (_row_5_d_x5_2_y),
    .z     (_row_5_d_x5_2_z)
  );
  ADD row_5_n_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:700:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_115_2092_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2110:118
    .y     (_row_5_d_x3_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:691:100
    .z     (_row_5_n_x7_2_z)
  );
  dup_2 row_5_d_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:701:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:700:100
    .y     (_row_5_d_x7_2_y),
    .z     (_row_5_d_x7_2_z)
  );
  SUB row_5_n_x8_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:702:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_115_2232_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2250:118
    .y     (_row_5_d_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:691:100
    .z     (_row_5_n_x8_4_z)
  );
  dup_2 row_5_d_x8_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:703:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x8_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:702:100
    .y     (_row_5_d_x8_4_y),
    .z     (_row_5_d_x8_4_z)
  );
  ADD row_5_n_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:704:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_141_2116_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2134:118
    .y     (_row_5_d_x2_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:688:100
    .z     (_row_5_n_x3_2_z)
  );
  dup_2 row_5_d_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:705:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:704:100
    .y     (_row_5_d_x3_2_y),
    .z     (_row_5_d_x3_2_z)
  );
  SUB row_5_n_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:706:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_141_2090_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2108:118
    .y     (_row_5_d_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:688:100
    .z     (_row_5_n_x0_2_z)
  );
  dup_2 row_5_d_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:707:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:706:100
    .y     (_row_5_d_x0_2_y),
    .z     (_row_5_d_x0_2_z)
  );
  ADD row_5_n_u2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:708:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_63_2089_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2107:114
    .y     (_row_5_d_x5_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:699:100
    .z     (_row_5_n_u2_2_z)
  );
  MUL row_5_n_v2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:709:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_c181_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:639:76
    .y     (_row_5_n_u2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:708:100
    .z     (_row_5_n_v2_2_z)
  );
  ADD row_5_n_w2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:710:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_v2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:709:100
    .y     (_row_5_n_c128_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:637:76
    .z     (_row_5_n_w2_2_z)
  );
  SHR_8 row_5_n_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:711:83
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_w2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:710:100
    .z     (_row_5_n_x2_2_z)
  );
  dup_2 row_5_d_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:712:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:711:83
    .y     (_row_5_d_x2_2_y),
    .z     (_row_5_d_x2_2_z)
  );
  SUB row_5_n_u4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:713:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_63_2190_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2208:114
    .y     (_row_5_d_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:699:100
    .z     (_row_5_n_u4_3_z)
  );
  MUL row_5_n_v4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:714:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_c181_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:640:76
    .y     (_row_5_n_u4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:713:100
    .z     (_row_5_n_v4_3_z)
  );
  ADD row_5_n_w4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:715:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_v4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:714:100
    .y     (_row_5_n_c128_2_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:638:76
    .z     (_row_5_n_w4_3_z)
  );
  SHR_8 row_5_n_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:716:83
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_w4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:715:100
    .z     (_row_5_n_x4_3_z)
  );
  dup_2 row_5_d_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:717:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:716:83
    .y     (_row_5_d_x4_3_y),
    .z     (_row_5_d_x4_3_z)
  );
  ADD row_5_n_tmp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:718:105
    .clock (clock),
    .reset (reset),
    .x     (_row_5_d_x7_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:701:100
    .y     (_delay_INT16_142_2088_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2106:118
    .z     (_row_5_n_tmp_0_z)
  );
  SHR_8 row_5_n_shr_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:719:87
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_tmp_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:718:105
    .z     (_row_5_n_shr_0_z)
  );
  ADD row_5_n_tmp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:720:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_134_2087_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2105:118
    .y     (_row_5_d_x2_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:712:100
    .z     (_row_5_n_tmp_1_z)
  );
  SHR_8 row_5_n_shr_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:721:87
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_tmp_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:720:105
    .z     (_row_5_n_shr_1_z)
  );
  ADD row_5_n_tmp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:722:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_134_2086_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2104:118
    .y     (_row_5_d_x4_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:717:100
    .z     (_row_5_n_tmp_2_z)
  );
  SHR_8 row_5_n_shr_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:723:87
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_tmp_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:722:105
    .z     (_row_5_n_shr_2_z)
  );
  ADD row_5_n_tmp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:724:105
    .clock (clock),
    .reset (reset),
    .x     (_row_5_d_x8_4_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:703:100
    .y     (_delay_INT16_184_2174_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2192:118
    .z     (_row_5_n_tmp_3_z)
  );
  SHR_8 row_5_n_shr_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:725:87
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_tmp_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:724:105
    .z     (_row_5_n_shr_3_z)
  );
  SUB row_5_n_tmp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:726:105
    .clock (clock),
    .reset (reset),
    .x     (_row_5_d_x8_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:703:100
    .y     (_delay_INT16_184_2185_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2203:118
    .z     (_row_5_n_tmp_4_z)
  );
  SHR_8 row_5_n_shr_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:727:87
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_tmp_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:726:105
    .z     (_row_5_n_shr_4_z)
  );
  SUB row_5_n_tmp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:728:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_134_2085_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2103:118
    .y     (_row_5_d_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:717:100
    .z     (_row_5_n_tmp_5_z)
  );
  SHR_8 row_5_n_shr_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:729:87
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_tmp_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:728:105
    .z     (_row_5_n_shr_5_z)
  );
  SUB row_5_n_tmp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:730:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_134_2084_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2102:118
    .y     (_row_5_d_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:712:100
    .z     (_row_5_n_tmp_6_z)
  );
  SHR_8 row_5_n_shr_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:731:87
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_tmp_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:730:105
    .z     (_row_5_n_shr_6_z)
  );
  SUB row_5_n_tmp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:732:105
    .clock (clock),
    .reset (reset),
    .x     (_row_5_d_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:701:100
    .y     (_delay_INT16_142_2306_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2324:118
    .z     (_row_5_n_tmp_7_z)
  );
  SHR_8 row_5_n_shr_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:733:87
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_tmp_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:732:105
    .z     (_row_5_n_shr_7_z)
  );
  C128 row_6_n_c128_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:734:76
    .clock (clock),
    .reset (reset),
    .value (_row_6_n_c128_0_value)
  );
  C128 row_6_n_c128_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:735:76
    .clock (clock),
    .reset (reset),
    .value (_row_6_n_c128_1_value)
  );
  C128 row_6_n_c128_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:736:76
    .clock (clock),
    .reset (reset),
    .value (_row_6_n_c128_2_value)
  );
  C181 row_6_n_c181_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:737:76
    .clock (clock),
    .reset (reset),
    .value (_row_6_n_c181_0_value)
  );
  C181 row_6_n_c181_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:738:76
    .clock (clock),
    .reset (reset),
    .value (_row_6_n_c181_1_value)
  );
  W7 row_6_n_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:739:64
    .clock (clock),
    .reset (reset),
    .value (_row_6_n_w7_value)
  );
  W1_sub_W7 row_6_n_w1_sub_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:740:85
    .clock (clock),
    .reset (reset),
    .value (_row_6_n_w1_sub_w7_value)
  );
  W1_add_W7 row_6_n_w1_add_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:741:85
    .clock (clock),
    .reset (reset),
    .value (_row_6_n_w1_add_w7_value)
  );
  W3 row_6_n_w3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:742:64
    .clock (clock),
    .reset (reset),
    .value (_row_6_n_w3_value)
  );
  W3_sub_W5 row_6_n_w3_sub_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:743:85
    .clock (clock),
    .reset (reset),
    .value (_row_6_n_w3_sub_w5_value)
  );
  W3_add_W5 row_6_n_w3_add_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:744:85
    .clock (clock),
    .reset (reset),
    .value (_row_6_n_w3_add_w5_value)
  );
  W6 row_6_n_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:745:64
    .clock (clock),
    .reset (reset),
    .value (_row_6_n_w6_value)
  );
  W2_sub_W6 row_6_n_w2_sub_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:746:85
    .clock (clock),
    .reset (reset),
    .value (_row_6_n_w2_sub_w6_value)
  );
  W2_add_W6 row_6_n_w2_add_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:747:85
    .clock (clock),
    .reset (reset),
    .value (_row_6_n_w2_add_w6_value)
  );
  SHL_11 row_6_n_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:748:83
    .clock (clock),
    .reset (reset),
    .x     (n_in_6_4_x),
    .z     (_row_6_n_x1_0_z)
  );
  SHL_11 row_6_n_t0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:749:83
    .clock (clock),
    .reset (reset),
    .x     (n_in_6_0_x),
    .z     (_row_6_n_t0_0_z)
  );
  ADD row_6_n_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:750:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_t0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:749:83
    .y     (_row_6_n_c128_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:734:76
    .z     (_row_6_n_x0_0_z)
  );
  dup_2 row_6_d_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:751:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:750:100
    .y     (_row_6_d_x0_0_y),
    .z     (_row_6_d_x0_0_z)
  );
  dup_2 row_6_d_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:752:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:748:83
    .y     (_row_6_d_x1_0_y),
    .z     (_row_6_d_x1_0_z)
  );
  dup_2 row_6_d_x2_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:753:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_6_6_x),
    .y     (_row_6_d_x2_0_y),
    .z     (_row_6_d_x2_0_z)
  );
  dup_2 row_6_d_x3_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:754:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_6_2_x),
    .y     (_row_6_d_x3_0_y),
    .z     (_row_6_d_x3_0_z)
  );
  dup_2 row_6_d_x4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:755:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_6_1_x),
    .y     (_row_6_d_x4_0_y),
    .z     (_row_6_d_x4_0_z)
  );
  dup_2 row_6_d_x5_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:756:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_6_7_x),
    .y     (_row_6_d_x5_0_y),
    .z     (_row_6_d_x5_0_z)
  );
  dup_2 row_6_d_x6_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:757:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_6_5_x),
    .y     (_row_6_d_x6_0_y),
    .z     (_row_6_d_x6_0_z)
  );
  dup_2 row_6_d_x7_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:758:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_6_3_x),
    .y     (_row_6_d_x7_0_y),
    .z     (_row_6_d_x7_0_z)
  );
  ADD row_6_n_t8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:759:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_47_2079_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2097:114
    .y     (_row_6_d_x5_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:756:100
    .z     (_row_6_n_t8_1_z)
  );
  MUL row_6_n_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:760:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:739:64
    .y     (_row_6_n_t8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:759:100
    .z     (_row_6_n_x8_1_z)
  );
  dup_2 row_6_d_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:761:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:760:100
    .y     (_row_6_d_x8_1_y),
    .z     (_row_6_d_x8_1_z)
  );
  MUL row_6_n_t4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:762:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_w1_sub_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:740:85
    .y     (_row_6_d_x4_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:755:100
    .z     (_row_6_n_t4_1_z)
  );
  ADD row_6_n_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:763:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_d_x8_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:761:100
    .y     (_delay_INT16_137_2278_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2296:118
    .z     (_row_6_n_x4_1_z)
  );
  dup_2 row_6_d_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:764:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:763:100
    .y     (_row_6_d_x4_1_y),
    .z     (_row_6_d_x4_1_z)
  );
  MUL row_6_n_t5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:765:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_w1_add_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:741:85
    .y     (_row_6_d_x5_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:756:100
    .z     (_row_6_n_t5_1_z)
  );
  SUB row_6_n_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:766:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_d_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:761:100
    .y     (_delay_INT16_173_2078_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2096:118
    .z     (_row_6_n_x5_1_z)
  );
  dup_2 row_6_d_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:767:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:766:100
    .y     (_row_6_d_x5_1_y),
    .z     (_row_6_d_x5_1_z)
  );
  ADD row_6_n_t8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:768:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_d_x6_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:757:100
    .y     (_delay_INT16_3_2077_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2095:110
    .z     (_row_6_n_t8_2_z)
  );
  MUL row_6_n_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:769:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_w3_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:742:64
    .y     (_row_6_n_t8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:768:100
    .z     (_row_6_n_x8_2_z)
  );
  dup_2 row_6_d_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:770:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:769:100
    .y     (_row_6_d_x8_2_y),
    .z     (_row_6_d_x8_2_z)
  );
  MUL row_6_n_t6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:771:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_w3_sub_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:743:85
    .y     (_row_6_d_x6_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:757:100
    .z     (_row_6_n_t6_1_z)
  );
  SUB row_6_n_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:772:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_d_x8_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:770:100
    .y     (_delay_INT16_139_2178_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2196:118
    .z     (_row_6_n_x6_1_z)
  );
  dup_2 row_6_d_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:773:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:772:100
    .y     (_row_6_d_x6_1_y),
    .z     (_row_6_d_x6_1_z)
  );
  MUL row_6_n_t7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:774:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_w3_add_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:744:85
    .y     (_row_6_d_x7_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:758:100
    .z     (_row_6_n_t7_1_z)
  );
  SUB row_6_n_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:775:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_d_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:770:100
    .y     (_delay_INT16_117_2127_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2145:118
    .z     (_row_6_n_x7_1_z)
  );
  dup_2 row_6_d_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:776:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:775:100
    .y     (_row_6_d_x7_1_y),
    .z     (_row_6_d_x7_1_z)
  );
  ADD row_6_n_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:777:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_d_x0_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:751:100
    .y     (_delay_INT16_39_2076_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2094:114
    .z     (_row_6_n_x8_3_z)
  );
  dup_2 row_6_d_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:778:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:777:100
    .y     (_row_6_d_x8_3_y),
    .z     (_row_6_d_x8_3_z)
  );
  SUB row_6_n_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:779:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_d_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:751:100
    .y     (_delay_INT16_39_2180_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2198:114
    .z     (_row_6_n_x0_1_z)
  );
  dup_2 row_6_d_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:780:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:779:100
    .y     (_row_6_d_x0_1_y),
    .z     (_row_6_d_x0_1_z)
  );
  ADD row_6_n_t1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:781:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_17_2075_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2093:114
    .y     (_row_6_d_x2_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:753:100
    .z     (_row_6_n_t1_1_z)
  );
  MUL row_6_n_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:782:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:745:64
    .y     (_row_6_n_t1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:781:100
    .z     (_row_6_n_x1_1_z)
  );
  dup_2 row_6_d_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:783:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:782:100
    .y     (_row_6_d_x1_1_y),
    .z     (_row_6_d_x1_1_z)
  );
  MUL row_6_n_t2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:784:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_w2_add_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:747:85
    .y     (_row_6_d_x2_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:753:100
    .z     (_row_6_n_t2_1_z)
  );
  SUB row_6_n_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:785:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_11_2074_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2092:114
    .y     (_row_6_n_t2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:784:100
    .z     (_row_6_n_x2_1_z)
  );
  dup_2 row_6_d_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:786:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:785:100
    .y     (_row_6_d_x2_1_y),
    .z     (_row_6_d_x2_1_z)
  );
  MUL row_6_n_t3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:787:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_w2_sub_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:746:85
    .y     (_row_6_d_x3_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:754:100
    .z     (_row_6_n_t3_1_z)
  );
  ADD row_6_n_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:788:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_26_2137_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2155:114
    .y     (_row_6_n_t3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:787:100
    .z     (_row_6_n_x3_1_z)
  );
  dup_2 row_6_d_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:789:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:788:100
    .y     (_row_6_d_x3_1_y),
    .z     (_row_6_d_x3_1_z)
  );
  ADD row_6_n_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:790:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_d_x4_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:764:100
    .y     (_delay_INT16_24_2072_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2090:114
    .z     (_row_6_n_x1_2_z)
  );
  dup_2 row_6_d_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:791:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:790:100
    .y     (_row_6_d_x1_2_y),
    .z     (_row_6_d_x1_2_z)
  );
  SUB row_6_n_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:792:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_d_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:764:100
    .y     (_delay_INT16_24_2071_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2089:114
    .z     (_row_6_n_x4_2_z)
  );
  dup_2 row_6_d_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:793:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:792:100
    .y     (_row_6_d_x4_2_y),
    .z     (_row_6_d_x4_2_z)
  );
  ADD row_6_n_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:794:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_d_x5_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:767:100
    .y     (_delay_INT16_17_2070_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2088:114
    .z     (_row_6_n_x6_2_z)
  );
  dup_2 row_6_d_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:795:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:794:100
    .y     (_row_6_d_x6_2_y),
    .z     (_row_6_d_x6_2_z)
  );
  SUB row_6_n_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:796:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_d_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:767:100
    .y     (_delay_INT16_17_2069_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2087:114
    .z     (_row_6_n_x5_2_z)
  );
  dup_2 row_6_d_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:797:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:796:100
    .y     (_row_6_d_x5_2_y),
    .z     (_row_6_d_x5_2_z)
  );
  ADD row_6_n_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:798:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_d_x8_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:778:100
    .y     (_delay_INT16_15_2068_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2086:114
    .z     (_row_6_n_x7_2_z)
  );
  dup_2 row_6_d_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:799:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:798:100
    .y     (_row_6_d_x7_2_y),
    .z     (_row_6_d_x7_2_z)
  );
  SUB row_6_n_x8_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:800:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_d_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:778:100
    .y     (_delay_INT16_15_2067_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2085:114
    .z     (_row_6_n_x8_4_z)
  );
  dup_2 row_6_d_x8_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:801:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x8_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:800:100
    .y     (_row_6_d_x8_4_y),
    .z     (_row_6_d_x8_4_z)
  );
  ADD row_6_n_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:802:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_d_x0_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:780:100
    .y     (_delay_INT16_14_2066_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2084:114
    .z     (_row_6_n_x3_2_z)
  );
  dup_2 row_6_d_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:803:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:802:100
    .y     (_row_6_d_x3_2_y),
    .z     (_row_6_d_x3_2_z)
  );
  SUB row_6_n_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:804:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_d_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:780:100
    .y     (_delay_INT16_14_2065_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2083:114
    .z     (_row_6_n_x0_2_z)
  );
  dup_2 row_6_d_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:805:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:804:100
    .y     (_row_6_d_x0_2_y),
    .z     (_row_6_d_x0_2_z)
  );
  ADD row_6_n_u2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:806:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_d_x4_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:793:100
    .y     (_delay_INT16_68_2064_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2082:114
    .z     (_row_6_n_u2_2_z)
  );
  MUL row_6_n_v2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:807:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_c181_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:737:76
    .y     (_row_6_n_u2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:806:100
    .z     (_row_6_n_v2_2_z)
  );
  ADD row_6_n_w2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:808:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_v2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:807:100
    .y     (_row_6_n_c128_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:735:76
    .z     (_row_6_n_w2_2_z)
  );
  SHR_8 row_6_n_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:809:83
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_w2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:808:100
    .z     (_row_6_n_x2_2_z)
  );
  dup_2 row_6_d_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:810:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:809:83
    .y     (_row_6_d_x2_2_y),
    .z     (_row_6_d_x2_2_z)
  );
  SUB row_6_n_u4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:811:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_d_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:793:100
    .y     (_delay_INT16_68_2133_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2151:114
    .z     (_row_6_n_u4_3_z)
  );
  MUL row_6_n_v4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:812:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_c181_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:738:76
    .y     (_row_6_n_u4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:811:100
    .z     (_row_6_n_v4_3_z)
  );
  ADD row_6_n_w4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:813:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_v4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:812:100
    .y     (_row_6_n_c128_2_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:736:76
    .z     (_row_6_n_w4_3_z)
  );
  SHR_8 row_6_n_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:814:83
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_w4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:813:100
    .z     (_row_6_n_x4_3_z)
  );
  dup_2 row_6_d_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:815:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:814:83
    .y     (_row_6_d_x4_3_y),
    .z     (_row_6_d_x4_3_z)
  );
  ADD row_6_n_tmp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:816:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_120_2063_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2081:118
    .y     (_row_6_d_x1_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:791:100
    .z     (_row_6_n_tmp_0_z)
  );
  SHR_8 row_6_n_shr_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:817:87
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_tmp_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:816:105
    .z     (_row_6_n_shr_0_z)
  );
  ADD row_6_n_tmp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:818:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_396_2062_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2080:118
    .y     (_row_6_d_x2_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:810:100
    .z     (_row_6_n_tmp_1_z)
  );
  SHR_8 row_6_n_shr_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:819:87
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_tmp_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:818:105
    .z     (_row_6_n_shr_1_z)
  );
  ADD row_6_n_tmp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:820:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_339_2142_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2160:118
    .y     (_row_6_d_x4_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:815:100
    .z     (_row_6_n_tmp_2_z)
  );
  SHR_8 row_6_n_shr_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:821:87
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_tmp_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:820:105
    .z     (_row_6_n_shr_2_z)
  );
  ADD row_6_n_tmp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:822:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_142_2061_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2079:118
    .y     (_row_6_d_x6_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:795:100
    .z     (_row_6_n_tmp_3_z)
  );
  SHR_8 row_6_n_shr_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:823:87
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_tmp_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:822:105
    .z     (_row_6_n_shr_3_z)
  );
  SUB row_6_n_tmp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:824:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_142_2060_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2078:118
    .y     (_row_6_d_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:795:100
    .z     (_row_6_n_tmp_4_z)
  );
  SHR_8 row_6_n_shr_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:825:87
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_tmp_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:824:105
    .z     (_row_6_n_shr_4_z)
  );
  SUB row_6_n_tmp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:826:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_339_2059_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2077:118
    .y     (_row_6_d_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:815:100
    .z     (_row_6_n_tmp_5_z)
  );
  SHR_8 row_6_n_shr_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:827:87
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_tmp_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:826:105
    .z     (_row_6_n_shr_5_z)
  );
  SUB row_6_n_tmp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:828:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_396_2057_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2075:118
    .y     (_row_6_d_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:810:100
    .z     (_row_6_n_tmp_6_z)
  );
  SHR_8 row_6_n_shr_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:829:87
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_tmp_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:828:105
    .z     (_row_6_n_shr_6_z)
  );
  SUB row_6_n_tmp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:830:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_120_2272_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2290:118
    .y     (_row_6_d_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:791:100
    .z     (_row_6_n_tmp_7_z)
  );
  SHR_8 row_6_n_shr_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:831:87
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_tmp_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:830:105
    .z     (_row_6_n_shr_7_z)
  );
  C128 row_7_n_c128_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:832:76
    .clock (clock),
    .reset (reset),
    .value (_row_7_n_c128_0_value)
  );
  C128 row_7_n_c128_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:833:76
    .clock (clock),
    .reset (reset),
    .value (_row_7_n_c128_1_value)
  );
  C128 row_7_n_c128_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:834:76
    .clock (clock),
    .reset (reset),
    .value (_row_7_n_c128_2_value)
  );
  C181 row_7_n_c181_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:835:76
    .clock (clock),
    .reset (reset),
    .value (_row_7_n_c181_0_value)
  );
  C181 row_7_n_c181_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:836:76
    .clock (clock),
    .reset (reset),
    .value (_row_7_n_c181_1_value)
  );
  W7 row_7_n_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:837:64
    .clock (clock),
    .reset (reset),
    .value (_row_7_n_w7_value)
  );
  W1_sub_W7 row_7_n_w1_sub_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:838:85
    .clock (clock),
    .reset (reset),
    .value (_row_7_n_w1_sub_w7_value)
  );
  W1_add_W7 row_7_n_w1_add_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:839:85
    .clock (clock),
    .reset (reset),
    .value (_row_7_n_w1_add_w7_value)
  );
  W3 row_7_n_w3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:840:64
    .clock (clock),
    .reset (reset),
    .value (_row_7_n_w3_value)
  );
  W3_sub_W5 row_7_n_w3_sub_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:841:85
    .clock (clock),
    .reset (reset),
    .value (_row_7_n_w3_sub_w5_value)
  );
  W3_add_W5 row_7_n_w3_add_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:842:85
    .clock (clock),
    .reset (reset),
    .value (_row_7_n_w3_add_w5_value)
  );
  W6 row_7_n_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:843:64
    .clock (clock),
    .reset (reset),
    .value (_row_7_n_w6_value)
  );
  W2_sub_W6 row_7_n_w2_sub_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:844:85
    .clock (clock),
    .reset (reset),
    .value (_row_7_n_w2_sub_w6_value)
  );
  W2_add_W6 row_7_n_w2_add_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:845:85
    .clock (clock),
    .reset (reset),
    .value (_row_7_n_w2_add_w6_value)
  );
  SHL_11 row_7_n_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:846:83
    .clock (clock),
    .reset (reset),
    .x     (n_in_7_4_x),
    .z     (_row_7_n_x1_0_z)
  );
  SHL_11 row_7_n_t0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:847:83
    .clock (clock),
    .reset (reset),
    .x     (n_in_7_0_x),
    .z     (_row_7_n_t0_0_z)
  );
  ADD row_7_n_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:848:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_t0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:847:83
    .y     (_row_7_n_c128_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:832:76
    .z     (_row_7_n_x0_0_z)
  );
  dup_2 row_7_d_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:849:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:848:100
    .y     (_row_7_d_x0_0_y),
    .z     (_row_7_d_x0_0_z)
  );
  dup_2 row_7_d_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:850:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:846:83
    .y     (_row_7_d_x1_0_y),
    .z     (_row_7_d_x1_0_z)
  );
  dup_2 row_7_d_x2_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:851:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_7_6_x),
    .y     (_row_7_d_x2_0_y),
    .z     (_row_7_d_x2_0_z)
  );
  dup_2 row_7_d_x3_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:852:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_7_2_x),
    .y     (_row_7_d_x3_0_y),
    .z     (_row_7_d_x3_0_z)
  );
  dup_2 row_7_d_x4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:853:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_7_1_x),
    .y     (_row_7_d_x4_0_y),
    .z     (_row_7_d_x4_0_z)
  );
  dup_2 row_7_d_x5_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:854:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_7_7_x),
    .y     (_row_7_d_x5_0_y),
    .z     (_row_7_d_x5_0_z)
  );
  dup_2 row_7_d_x6_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:855:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_7_5_x),
    .y     (_row_7_d_x6_0_y),
    .z     (_row_7_d_x6_0_z)
  );
  dup_2 row_7_d_x7_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:856:100
    .clock (clock),
    .reset (reset),
    .x     (n_in_7_3_x),
    .y     (_row_7_d_x7_0_y),
    .z     (_row_7_d_x7_0_z)
  );
  ADD row_7_n_t8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:857:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_d_x4_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:853:100
    .y     (_delay_INT16_19_2055_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2073:114
    .z     (_row_7_n_t8_1_z)
  );
  MUL row_7_n_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:858:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:837:64
    .y     (_row_7_n_t8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:857:100
    .z     (_row_7_n_x8_1_z)
  );
  dup_2 row_7_d_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:859:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:858:100
    .y     (_row_7_d_x8_1_y),
    .z     (_row_7_d_x8_1_z)
  );
  MUL row_7_n_t4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:860:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_w1_sub_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:838:85
    .y     (_row_7_d_x4_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:853:100
    .z     (_row_7_n_t4_1_z)
  );
  ADD row_7_n_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:861:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_d_x8_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:859:100
    .y     (_delay_INT16_34_2053_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2071:114
    .z     (_row_7_n_x4_1_z)
  );
  dup_2 row_7_d_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:862:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:861:100
    .y     (_row_7_d_x4_1_y),
    .z     (_row_7_d_x4_1_z)
  );
  MUL row_7_n_t5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:863:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_w1_add_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:839:85
    .y     (_row_7_d_x5_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:854:100
    .z     (_row_7_n_t5_1_z)
  );
  SUB row_7_n_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:864:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_d_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:859:100
    .y     (_delay_INT16_111_2050_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2068:118
    .z     (_row_7_n_x5_1_z)
  );
  dup_2 row_7_d_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:865:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:864:100
    .y     (_row_7_d_x5_1_y),
    .z     (_row_7_d_x5_1_z)
  );
  ADD row_7_n_t8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:866:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_d_x6_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:855:100
    .y     (_delay_INT16_1_2049_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2067:110
    .z     (_row_7_n_t8_2_z)
  );
  MUL row_7_n_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:867:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_w3_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:840:64
    .y     (_row_7_n_t8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:866:100
    .z     (_row_7_n_x8_2_z)
  );
  dup_2 row_7_d_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:868:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:867:100
    .y     (_row_7_d_x8_2_y),
    .z     (_row_7_d_x8_2_z)
  );
  MUL row_7_n_t6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:869:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_w3_sub_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:841:85
    .y     (_row_7_d_x6_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:855:100
    .z     (_row_7_n_t6_1_z)
  );
  SUB row_7_n_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:870:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_d_x8_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:868:100
    .y     (_delay_INT16_182_2047_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2065:118
    .z     (_row_7_n_x6_1_z)
  );
  dup_2 row_7_d_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:871:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:870:100
    .y     (_row_7_d_x6_1_y),
    .z     (_row_7_d_x6_1_z)
  );
  MUL row_7_n_t7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:872:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_w3_add_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:842:85
    .y     (_row_7_d_x7_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:856:100
    .z     (_row_7_n_t7_1_z)
  );
  SUB row_7_n_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:873:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_d_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:868:100
    .y     (_delay_INT16_147_2046_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2064:118
    .z     (_row_7_n_x7_1_z)
  );
  dup_2 row_7_d_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:874:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:873:100
    .y     (_row_7_d_x7_1_y),
    .z     (_row_7_d_x7_1_z)
  );
  ADD row_7_n_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:875:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_48_2146_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2164:114
    .y     (_row_7_d_x1_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:850:100
    .z     (_row_7_n_x8_3_z)
  );
  dup_2 row_7_d_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:876:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:875:100
    .y     (_row_7_d_x8_3_y),
    .z     (_row_7_d_x8_3_z)
  );
  SUB row_7_n_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:877:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_48_2044_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2062:114
    .y     (_row_7_d_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:850:100
    .z     (_row_7_n_x0_1_z)
  );
  dup_2 row_7_d_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:878:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:877:100
    .y     (_row_7_d_x0_1_y),
    .z     (_row_7_d_x0_1_z)
  );
  ADD row_7_n_t1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:879:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_d_x3_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:852:100
    .y     (_delay_INT16_121_2043_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2061:118
    .z     (_row_7_n_t1_1_z)
  );
  MUL row_7_n_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:880:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:843:64
    .y     (_row_7_n_t1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:879:100
    .z     (_row_7_n_x1_1_z)
  );
  dup_2 row_7_d_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:881:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:880:100
    .y     (_row_7_d_x1_1_y),
    .z     (_row_7_d_x1_1_z)
  );
  MUL row_7_n_t2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:882:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_w2_add_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:845:85
    .y     (_delay_INT16_13_2041_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2059:114
    .z     (_row_7_n_t2_1_z)
  );
  SUB row_7_n_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:883:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_d_x1_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:881:100
    .y     (_delay_INT16_100_2040_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2058:118
    .z     (_row_7_n_x2_1_z)
  );
  dup_2 row_7_d_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:884:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:883:100
    .y     (_row_7_d_x2_1_y),
    .z     (_row_7_d_x2_1_z)
  );
  MUL row_7_n_t3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:885:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_w2_sub_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:844:85
    .y     (_row_7_d_x3_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:852:100
    .z     (_row_7_n_t3_1_z)
  );
  ADD row_7_n_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:886:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_2_2302_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2320:110
    .y     (_row_7_n_t3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:885:100
    .z     (_row_7_n_x3_1_z)
  );
  dup_2 row_7_d_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:887:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:886:100
    .y     (_row_7_d_x3_1_y),
    .z     (_row_7_d_x3_1_z)
  );
  ADD row_7_n_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:888:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_33_2039_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2057:114
    .y     (_row_7_d_x6_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:871:100
    .z     (_row_7_n_x1_2_z)
  );
  dup_2 row_7_d_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:889:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:888:100
    .y     (_row_7_d_x1_2_y),
    .z     (_row_7_d_x1_2_z)
  );
  SUB row_7_n_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:890:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_33_2093_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2111:114
    .y     (_row_7_d_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:871:100
    .z     (_row_7_n_x4_2_z)
  );
  dup_2 row_7_d_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:891:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:890:100
    .y     (_row_7_d_x4_2_y),
    .z     (_row_7_d_x4_2_z)
  );
  ADD row_7_n_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:892:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_35_2038_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2056:114
    .y     (_row_7_d_x7_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:874:100
    .z     (_row_7_n_x6_2_z)
  );
  dup_2 row_7_d_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:893:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:892:100
    .y     (_row_7_d_x6_2_y),
    .z     (_row_7_d_x6_2_z)
  );
  SUB row_7_n_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:894:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_35_2037_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2055:114
    .y     (_row_7_d_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:874:100
    .z     (_row_7_n_x5_2_z)
  );
  dup_2 row_7_d_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:895:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:894:100
    .y     (_row_7_d_x5_2_y),
    .z     (_row_7_d_x5_2_z)
  );
  ADD row_7_n_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:896:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_d_x8_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:876:100
    .y     (_delay_INT16_6_2251_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2269:110
    .z     (_row_7_n_x7_2_z)
  );
  dup_2 row_7_d_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:897:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:896:100
    .y     (_row_7_d_x7_2_y),
    .z     (_row_7_d_x7_2_z)
  );
  SUB row_7_n_x8_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:898:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_d_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:876:100
    .y     (_delay_INT16_6_2036_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2054:110
    .z     (_row_7_n_x8_4_z)
  );
  dup_2 row_7_d_x8_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:899:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x8_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:898:100
    .y     (_row_7_d_x8_4_y),
    .z     (_row_7_d_x8_4_z)
  );
  ADD row_7_n_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:900:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_19_2035_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2053:114
    .y     (_row_7_d_x2_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:884:100
    .z     (_row_7_n_x3_2_z)
  );
  dup_2 row_7_d_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:901:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:900:100
    .y     (_row_7_d_x3_2_y),
    .z     (_row_7_d_x3_2_z)
  );
  SUB row_7_n_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:902:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_19_2316_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2334:114
    .y     (_row_7_d_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:884:100
    .z     (_row_7_n_x0_2_z)
  );
  dup_2 row_7_d_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:903:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:902:100
    .y     (_row_7_d_x0_2_y),
    .z     (_row_7_d_x0_2_z)
  );
  ADD row_7_n_u2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:904:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_d_x4_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:891:100
    .y     (_delay_INT16_13_2033_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2051:114
    .z     (_row_7_n_u2_2_z)
  );
  MUL row_7_n_v2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:905:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_c181_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:835:76
    .y     (_row_7_n_u2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:904:100
    .z     (_row_7_n_v2_2_z)
  );
  ADD row_7_n_w2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:906:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_v2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:905:100
    .y     (_row_7_n_c128_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:833:76
    .z     (_row_7_n_w2_2_z)
  );
  SHR_8 row_7_n_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:907:83
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_w2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:906:100
    .z     (_row_7_n_x2_2_z)
  );
  dup_2 row_7_d_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:908:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:907:83
    .y     (_row_7_d_x2_2_y),
    .z     (_row_7_d_x2_2_z)
  );
  SUB row_7_n_u4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:909:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_d_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:891:100
    .y     (_delay_INT16_13_2032_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2050:114
    .z     (_row_7_n_u4_3_z)
  );
  MUL row_7_n_v4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:910:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_c181_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:836:76
    .y     (_row_7_n_u4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:909:100
    .z     (_row_7_n_v4_3_z)
  );
  ADD row_7_n_w4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:911:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_v4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:910:100
    .y     (_row_7_n_c128_2_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:834:76
    .z     (_row_7_n_w4_3_z)
  );
  SHR_8 row_7_n_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:912:83
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_w4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:911:100
    .z     (_row_7_n_x4_3_z)
  );
  dup_2 row_7_d_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:913:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:912:83
    .y     (_row_7_d_x4_3_y),
    .z     (_row_7_d_x4_3_z)
  );
  ADD row_7_n_tmp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:914:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_45_2031_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2049:114
    .y     (_row_7_d_x1_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:889:100
    .z     (_row_7_n_tmp_0_z)
  );
  SHR_8 row_7_n_shr_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:915:87
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_tmp_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:914:105
    .z     (_row_7_n_shr_0_z)
  );
  ADD row_7_n_tmp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:916:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_338_2030_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2048:118
    .y     (_row_7_d_x2_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:908:100
    .z     (_row_7_n_tmp_1_z)
  );
  SHR_8 row_7_n_shr_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:917:87
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_tmp_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:916:105
    .z     (_row_7_n_shr_1_z)
  );
  ADD row_7_n_tmp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:918:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_255_2029_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2047:118
    .y     (_row_7_d_x4_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:913:100
    .z     (_row_7_n_tmp_2_z)
  );
  SHR_8 row_7_n_shr_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:919:87
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_tmp_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:918:105
    .z     (_row_7_n_shr_2_z)
  );
  ADD row_7_n_tmp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:920:105
    .clock (clock),
    .reset (reset),
    .x     (_row_7_d_x8_4_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:899:100
    .y     (_delay_INT16_122_2028_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2046:118
    .z     (_row_7_n_tmp_3_z)
  );
  SHR_8 row_7_n_shr_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:921:87
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_tmp_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:920:105
    .z     (_row_7_n_shr_3_z)
  );
  SUB row_7_n_tmp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:922:105
    .clock (clock),
    .reset (reset),
    .x     (_row_7_d_x8_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:899:100
    .y     (_delay_INT16_122_2027_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2045:118
    .z     (_row_7_n_tmp_4_z)
  );
  SHR_8 row_7_n_shr_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:923:87
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_tmp_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:922:105
    .z     (_row_7_n_shr_4_z)
  );
  SUB row_7_n_tmp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:924:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_255_2026_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2044:118
    .y     (_row_7_d_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:913:100
    .z     (_row_7_n_tmp_5_z)
  );
  SHR_8 row_7_n_shr_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:925:87
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_tmp_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:924:105
    .z     (_row_7_n_shr_5_z)
  );
  SUB row_7_n_tmp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:926:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_338_2024_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2042:118
    .y     (_row_7_d_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:908:100
    .z     (_row_7_n_tmp_6_z)
  );
  SHR_8 row_7_n_shr_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:927:87
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_tmp_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:926:105
    .z     (_row_7_n_shr_6_z)
  );
  SUB row_7_n_tmp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:928:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_45_2023_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2041:114
    .y     (_row_7_d_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:889:100
    .z     (_row_7_n_tmp_7_z)
  );
  SHR_8 row_7_n_shr_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:929:87
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_tmp_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:928:105
    .z     (_row_7_n_shr_7_z)
  );
  C4 col_0_n_c4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:930:70
    .clock (clock),
    .reset (reset),
    .value (_col_0_n_c4_0_value)
  );
  C4 col_0_n_c4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:931:70
    .clock (clock),
    .reset (reset),
    .value (_col_0_n_c4_1_value)
  );
  C4 col_0_n_c4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:932:70
    .clock (clock),
    .reset (reset),
    .value (_col_0_n_c4_2_value)
  );
  C128 col_0_n_c128_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:933:76
    .clock (clock),
    .reset (reset),
    .value (_col_0_n_c128_0_value)
  );
  C128 col_0_n_c128_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:934:76
    .clock (clock),
    .reset (reset),
    .value (_col_0_n_c128_1_value)
  );
  C181 col_0_n_c181_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:935:76
    .clock (clock),
    .reset (reset),
    .value (_col_0_n_c181_0_value)
  );
  C181 col_0_n_c181_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:936:76
    .clock (clock),
    .reset (reset),
    .value (_col_0_n_c181_1_value)
  );
  C8192 col_0_n_c8192 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:937:73
    .clock (clock),
    .reset (reset),
    .value (_col_0_n_c8192_value)
  );
  W7 col_0_n_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:938:64
    .clock (clock),
    .reset (reset),
    .value (_col_0_n_w7_value)
  );
  W1_sub_W7 col_0_n_w1_sub_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:939:85
    .clock (clock),
    .reset (reset),
    .value (_col_0_n_w1_sub_w7_value)
  );
  W1_add_W7 col_0_n_w1_add_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:940:85
    .clock (clock),
    .reset (reset),
    .value (_col_0_n_w1_add_w7_value)
  );
  W3 col_0_n_w3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:941:64
    .clock (clock),
    .reset (reset),
    .value (_col_0_n_w3_value)
  );
  W3_sub_W5 col_0_n_w3_sub_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:942:85
    .clock (clock),
    .reset (reset),
    .value (_col_0_n_w3_sub_w5_value)
  );
  W3_add_W5 col_0_n_w3_add_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:943:85
    .clock (clock),
    .reset (reset),
    .value (_col_0_n_w3_add_w5_value)
  );
  W6 col_0_n_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:944:64
    .clock (clock),
    .reset (reset),
    .value (_col_0_n_w6_value)
  );
  W2_sub_W6 col_0_n_w2_sub_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:945:85
    .clock (clock),
    .reset (reset),
    .value (_col_0_n_w2_sub_w6_value)
  );
  W2_add_W6 col_0_n_w2_add_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:946:85
    .clock (clock),
    .reset (reset),
    .value (_col_0_n_w2_add_w6_value)
  );
  SHL_8 col_0_n_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:947:83
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_shr_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:621:87
    .z     (_col_0_n_x1_0_z)
  );
  SHL_8 col_0_n_t0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:948:83
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_shr_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:229:87
    .z     (_col_0_n_t0_0_z)
  );
  ADD col_0_n_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:949:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_t0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:948:83
    .y     (_col_0_n_c8192_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:937:73
    .z     (_col_0_n_x0_0_z)
  );
  dup_2 col_0_d_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:950:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:949:100
    .y     (_col_0_d_x0_0_y),
    .z     (_col_0_d_x0_0_z)
  );
  dup_2 col_0_d_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:951:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:947:83
    .y     (_col_0_d_x1_0_y),
    .z     (_col_0_d_x1_0_z)
  );
  dup_2 col_0_d_x2_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:952:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_shr_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:817:87
    .y     (_col_0_d_x2_0_y),
    .z     (_col_0_d_x2_0_z)
  );
  dup_2 col_0_d_x3_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:953:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_shr_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:425:87
    .y     (_col_0_d_x3_0_y),
    .z     (_col_0_d_x3_0_z)
  );
  dup_2 col_0_d_x4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:954:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_shr_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:327:87
    .y     (_col_0_d_x4_0_y),
    .z     (_col_0_d_x4_0_z)
  );
  dup_2 col_0_d_x5_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:955:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_shr_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:915:87
    .y     (_col_0_d_x5_0_y),
    .z     (_col_0_d_x5_0_z)
  );
  dup_2 col_0_d_x6_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:956:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_shr_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:719:87
    .y     (_col_0_d_x6_0_y),
    .z     (_col_0_d_x6_0_z)
  );
  dup_2 col_0_d_x7_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:957:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_shr_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:523:87
    .y     (_col_0_d_x7_0_y),
    .z     (_col_0_d_x7_0_z)
  );
  ADD col_0_n_u8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:958:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_7_2019_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2037:110
    .y     (_col_0_d_x5_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:955:100
    .z     (_col_0_n_u8_0_z)
  );
  MUL col_0_n_v8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:959:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:938:64
    .y     (_col_0_n_u8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:958:100
    .z     (_col_0_n_v8_0_z)
  );
  ADD col_0_n_x8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:960:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_v8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:959:100
    .y     (_col_0_n_c4_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:930:70
    .z     (_col_0_n_x8_0_z)
  );
  dup_2 col_0_d_x8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:961:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:960:100
    .y     (_col_0_d_x8_0_y),
    .z     (_col_0_d_x8_0_z)
  );
  MUL col_0_n_u4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:962:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_w1_sub_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:939:85
    .y     (_col_0_d_x4_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:954:100
    .z     (_col_0_n_u4_1_z)
  );
  ADD col_0_n_v4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:963:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_d_x8_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:961:100
    .y     (_delay_INT16_217_2209_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2227:118
    .z     (_col_0_n_v4_1_z)
  );
  SHR_3 col_0_n_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:964:83
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_v4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:963:100
    .z     (_col_0_n_x4_1_z)
  );
  dup_2 col_0_d_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:965:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:964:83
    .y     (_col_0_d_x4_1_y),
    .z     (_col_0_d_x4_1_z)
  );
  MUL col_0_n_u5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:966:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_w1_add_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:940:85
    .y     (_col_0_d_x5_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:955:100
    .z     (_col_0_n_u5_1_z)
  );
  SUB col_0_n_v5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:967:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_d_x8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:961:100
    .y     (_delay_INT16_298_2017_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2035:118
    .z     (_col_0_n_v5_1_z)
  );
  SHR_3 col_0_n_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:968:83
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_v5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:967:100
    .z     (_col_0_n_x5_1_z)
  );
  dup_2 col_0_d_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:969:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:968:83
    .y     (_col_0_d_x5_1_y),
    .z     (_col_0_d_x5_1_z)
  );
  ADD col_0_n_u8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:970:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_181_2016_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2034:118
    .y     (_col_0_d_x7_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:957:100
    .z     (_col_0_n_u8_1_z)
  );
  MUL col_0_n_v8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:971:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_w3_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:941:64
    .y     (_col_0_n_u8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:970:100
    .z     (_col_0_n_v8_1_z)
  );
  ADD col_0_n_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:972:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_v8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:971:100
    .y     (_col_0_n_c4_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:931:70
    .z     (_col_0_n_x8_1_z)
  );
  dup_2 col_0_d_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:973:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:972:100
    .y     (_col_0_d_x8_1_y),
    .z     (_col_0_d_x8_1_z)
  );
  MUL col_0_n_u6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:974:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_w3_sub_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:942:85
    .y     (_col_0_d_x6_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:956:100
    .z     (_col_0_n_u6_1_z)
  );
  SUB col_0_n_v6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:975:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_d_x8_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:973:100
    .y     (_delay_INT16_370_2123_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2141:118
    .z     (_col_0_n_v6_1_z)
  );
  SHR_3 col_0_n_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:976:83
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_v6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:975:100
    .z     (_col_0_n_x6_1_z)
  );
  dup_2 col_0_d_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:977:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:976:83
    .y     (_col_0_d_x6_1_y),
    .z     (_col_0_d_x6_1_z)
  );
  MUL col_0_n_u7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:978:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_w3_add_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:943:85
    .y     (_col_0_d_x7_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:957:100
    .z     (_col_0_n_u7_1_z)
  );
  SUB col_0_n_v7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:979:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_d_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:973:100
    .y     (_delay_INT16_185_2135_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2153:118
    .z     (_col_0_n_v7_1_z)
  );
  SHR_3 col_0_n_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:980:83
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_v7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:979:100
    .z     (_col_0_n_x7_1_z)
  );
  dup_2 col_0_d_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:981:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:980:83
    .y     (_col_0_d_x7_1_y),
    .z     (_col_0_d_x7_1_z)
  );
  ADD col_0_n_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:982:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_242_2014_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2032:118
    .y     (_col_0_d_x1_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:951:100
    .z     (_col_0_n_x8_2_z)
  );
  dup_2 col_0_d_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:983:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:982:100
    .y     (_col_0_d_x8_2_y),
    .z     (_col_0_d_x8_2_z)
  );
  SUB col_0_n_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:984:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_242_2012_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2030:118
    .y     (_col_0_d_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:951:100
    .z     (_col_0_n_x0_1_z)
  );
  dup_2 col_0_d_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:985:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:984:100
    .y     (_col_0_d_x0_1_y),
    .z     (_col_0_d_x0_1_z)
  );
  ADD col_0_n_u1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:986:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_158_2311_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2329:118
    .y     (_col_0_d_x2_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:952:100
    .z     (_col_0_n_u1_1_z)
  );
  MUL col_0_n_v1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:987:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:944:64
    .y     (_col_0_n_u1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:986:100
    .z     (_col_0_n_v1_1_z)
  );
  ADD col_0_n_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:988:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_v1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:987:100
    .y     (_col_0_n_c4_2_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:932:70
    .z     (_col_0_n_x1_1_z)
  );
  dup_2 col_0_d_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:989:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:988:100
    .y     (_col_0_d_x1_1_y),
    .z     (_col_0_d_x1_1_z)
  );
  MUL col_0_n_u2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:990:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_w2_add_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:946:85
    .y     (_col_0_d_x2_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:952:100
    .z     (_col_0_n_u2_1_z)
  );
  SUB col_0_n_v2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:991:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_d_x1_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:989:100
    .y     (_delay_INT16_127_2011_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2029:118
    .z     (_col_0_n_v2_1_z)
  );
  SHR_3 col_0_n_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:992:83
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_v2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:991:100
    .z     (_col_0_n_x2_1_z)
  );
  dup_2 col_0_d_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:993:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:992:83
    .y     (_col_0_d_x2_1_y),
    .z     (_col_0_d_x2_1_z)
  );
  MUL col_0_n_u3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:994:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_w2_sub_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:945:85
    .y     (_col_0_d_x3_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:953:100
    .z     (_col_0_n_u3_1_z)
  );
  ADD col_0_n_v3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:995:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_d_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:989:100
    .y     (_delay_INT16_296_2009_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2027:118
    .z     (_col_0_n_v3_1_z)
  );
  SHR_3 col_0_n_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:996:83
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_v3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:995:100
    .z     (_col_0_n_x3_1_z)
  );
  dup_2 col_0_d_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:997:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:996:83
    .y     (_col_0_d_x3_1_y),
    .z     (_col_0_d_x3_1_z)
  );
  ADD col_0_n_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:998:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_212_2007_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2025:118
    .y     (_col_0_d_x6_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:977:100
    .z     (_col_0_n_x1_2_z)
  );
  dup_2 col_0_d_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:999:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:998:100
    .y     (_col_0_d_x1_2_y),
    .z     (_col_0_d_x1_2_z)
  );
  SUB col_0_n_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1000:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_212_2006_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2024:118
    .y     (_col_0_d_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:977:100
    .z     (_col_0_n_x4_2_z)
  );
  dup_2 col_0_d_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1001:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1000:100
    .y     (_col_0_d_x4_2_y),
    .z     (_col_0_d_x4_2_z)
  );
  ADD col_0_n_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1002:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_94_2004_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2022:114
    .y     (_col_0_d_x7_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:981:100
    .z     (_col_0_n_x6_2_z)
  );
  dup_2 col_0_d_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1003:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1002:100
    .y     (_col_0_d_x6_2_y),
    .z     (_col_0_d_x6_2_z)
  );
  SUB col_0_n_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1004:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_94_2002_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2020:114
    .y     (_col_0_d_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:981:100
    .z     (_col_0_n_x5_2_z)
  );
  dup_2 col_0_d_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1005:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1004:100
    .y     (_col_0_d_x5_2_y),
    .z     (_col_0_d_x5_2_z)
  );
  ADD col_0_n_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1006:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_139_2001_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2019:118
    .y     (_col_0_d_x3_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:997:100
    .z     (_col_0_n_x7_2_z)
  );
  dup_2 col_0_d_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1007:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1006:100
    .y     (_col_0_d_x7_2_y),
    .z     (_col_0_d_x7_2_z)
  );
  SUB col_0_n_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1008:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_139_2000_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2018:118
    .y     (_col_0_d_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:997:100
    .z     (_col_0_n_x8_3_z)
  );
  dup_2 col_0_d_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1009:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1008:100
    .y     (_col_0_d_x8_3_y),
    .z     (_col_0_d_x8_3_z)
  );
  ADD col_0_n_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1010:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_23_1999_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2017:114
    .y     (_col_0_d_x2_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:993:100
    .z     (_col_0_n_x3_2_z)
  );
  dup_2 col_0_d_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1011:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1010:100
    .y     (_col_0_d_x3_2_y),
    .z     (_col_0_d_x3_2_z)
  );
  SUB col_0_n_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1012:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_23_1998_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2016:114
    .y     (_col_0_d_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:993:100
    .z     (_col_0_n_x0_2_z)
  );
  dup_2 col_0_d_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1013:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1012:100
    .y     (_col_0_d_x0_2_y),
    .z     (_col_0_d_x0_2_z)
  );
  ADD col_0_n_u2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1014:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_d_x4_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1001:100
    .y     (_delay_INT16_89_1997_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2015:114
    .z     (_col_0_n_u2_2_z)
  );
  MUL col_0_n_v2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1015:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_c181_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:935:76
    .y     (_col_0_n_u2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1014:100
    .z     (_col_0_n_v2_2_z)
  );
  ADD col_0_n_w2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1016:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_v2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1015:100
    .y     (_col_0_n_c128_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:933:76
    .z     (_col_0_n_w2_2_z)
  );
  SHR_8 col_0_n_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1017:83
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_w2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1016:100
    .z     (_col_0_n_x2_2_z)
  );
  dup_2 col_0_d_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1018:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1017:83
    .y     (_col_0_d_x2_2_y),
    .z     (_col_0_d_x2_2_z)
  );
  SUB col_0_n_u4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1019:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_d_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1001:100
    .y     (_delay_INT16_89_1996_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2014:114
    .z     (_col_0_n_u4_3_z)
  );
  MUL col_0_n_v4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1020:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_c181_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:936:76
    .y     (_col_0_n_u4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1019:100
    .z     (_col_0_n_v4_3_z)
  );
  ADD col_0_n_w4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1021:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_v4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1020:100
    .y     (_col_0_n_c128_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:934:76
    .z     (_col_0_n_w4_3_z)
  );
  SHR_8 col_0_n_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1022:83
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_w4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1021:100
    .z     (_col_0_n_x4_3_z)
  );
  dup_2 col_0_d_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1023:100
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1022:83
    .y     (_col_0_d_x4_3_y),
    .z     (_col_0_d_x4_3_z)
  );
  ADD col_0_n_tmp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1024:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_94_1995_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2013:114
    .y     (_col_0_d_x1_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:999:100
    .z     (_col_0_n_tmp_0_z)
  );
  SHR_14 col_0_n_val_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1025:87
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_tmp_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1024:105
    .z     (_col_0_n_val_0_z)
  );
  CLIP col_0_n_clp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1026:87
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_val_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1025:87
    .z     (n_out_0_0_x)
  );
  ADD col_0_n_tmp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1027:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_487_1994_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2012:118
    .y     (_col_0_d_x2_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1018:100
    .z     (_col_0_n_tmp_1_z)
  );
  SHR_14 col_0_n_val_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1028:87
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_tmp_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1027:105
    .z     (_col_0_n_val_1_z)
  );
  CLIP col_0_n_clp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1029:87
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_val_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1028:87
    .z     (n_out_1_0_x)
  );
  ADD col_0_n_tmp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1030:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_477_2151_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2169:118
    .y     (_col_0_d_x4_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1023:100
    .z     (_col_0_n_tmp_2_z)
  );
  SHR_14 col_0_n_val_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1031:87
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_tmp_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1030:105
    .z     (_col_0_n_val_2_z)
  );
  CLIP col_0_n_clp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1032:87
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_val_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1031:87
    .z     (n_out_2_0_x)
  );
  ADD col_0_n_tmp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1033:105
    .clock (clock),
    .reset (reset),
    .x     (_col_0_d_x8_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1009:100
    .y     (_delay_INT16_34_1993_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2011:114
    .z     (_col_0_n_tmp_3_z)
  );
  SHR_14 col_0_n_val_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1034:87
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_tmp_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1033:105
    .z     (_col_0_n_val_3_z)
  );
  CLIP col_0_n_clp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1035:87
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_val_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1034:87
    .z     (n_out_3_0_x)
  );
  SUB col_0_n_tmp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1036:105
    .clock (clock),
    .reset (reset),
    .x     (_col_0_d_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1009:100
    .y     (_delay_INT16_34_2315_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2333:114
    .z     (_col_0_n_tmp_4_z)
  );
  SHR_14 col_0_n_val_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1037:87
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_tmp_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1036:105
    .z     (_col_0_n_val_4_z)
  );
  CLIP col_0_n_clp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1038:87
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_val_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1037:87
    .z     (n_out_4_0_x)
  );
  SUB col_0_n_tmp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1039:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_477_1992_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2010:118
    .y     (_col_0_d_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1023:100
    .z     (_col_0_n_tmp_5_z)
  );
  SHR_14 col_0_n_val_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1040:87
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_tmp_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1039:105
    .z     (_col_0_n_val_5_z)
  );
  CLIP col_0_n_clp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1041:87
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_val_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1040:87
    .z     (n_out_5_0_x)
  );
  SUB col_0_n_tmp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1042:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_487_1991_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2009:118
    .y     (_col_0_d_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1018:100
    .z     (_col_0_n_tmp_6_z)
  );
  SHR_14 col_0_n_val_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1043:87
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_tmp_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1042:105
    .z     (_col_0_n_val_6_z)
  );
  CLIP col_0_n_clp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1044:87
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_val_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1043:87
    .z     (n_out_6_0_x)
  );
  SUB col_0_n_tmp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1045:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_94_1990_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2008:114
    .y     (_col_0_d_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:999:100
    .z     (_col_0_n_tmp_7_z)
  );
  SHR_14 col_0_n_val_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1046:87
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_tmp_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1045:105
    .z     (_col_0_n_val_7_z)
  );
  CLIP col_0_n_clp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1047:87
    .clock (clock),
    .reset (reset),
    .x     (_col_0_n_val_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1046:87
    .z     (n_out_7_0_x)
  );
  C4 col_1_n_c4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1048:70
    .clock (clock),
    .reset (reset),
    .value (_col_1_n_c4_0_value)
  );
  C4 col_1_n_c4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1049:70
    .clock (clock),
    .reset (reset),
    .value (_col_1_n_c4_1_value)
  );
  C4 col_1_n_c4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1050:70
    .clock (clock),
    .reset (reset),
    .value (_col_1_n_c4_2_value)
  );
  C128 col_1_n_c128_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1051:76
    .clock (clock),
    .reset (reset),
    .value (_col_1_n_c128_0_value)
  );
  C128 col_1_n_c128_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1052:76
    .clock (clock),
    .reset (reset),
    .value (_col_1_n_c128_1_value)
  );
  C181 col_1_n_c181_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1053:76
    .clock (clock),
    .reset (reset),
    .value (_col_1_n_c181_0_value)
  );
  C181 col_1_n_c181_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1054:76
    .clock (clock),
    .reset (reset),
    .value (_col_1_n_c181_1_value)
  );
  C8192 col_1_n_c8192 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1055:73
    .clock (clock),
    .reset (reset),
    .value (_col_1_n_c8192_value)
  );
  W7 col_1_n_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1056:64
    .clock (clock),
    .reset (reset),
    .value (_col_1_n_w7_value)
  );
  W1_sub_W7 col_1_n_w1_sub_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1057:85
    .clock (clock),
    .reset (reset),
    .value (_col_1_n_w1_sub_w7_value)
  );
  W1_add_W7 col_1_n_w1_add_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1058:85
    .clock (clock),
    .reset (reset),
    .value (_col_1_n_w1_add_w7_value)
  );
  W3 col_1_n_w3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1059:64
    .clock (clock),
    .reset (reset),
    .value (_col_1_n_w3_value)
  );
  W3_sub_W5 col_1_n_w3_sub_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1060:85
    .clock (clock),
    .reset (reset),
    .value (_col_1_n_w3_sub_w5_value)
  );
  W3_add_W5 col_1_n_w3_add_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1061:85
    .clock (clock),
    .reset (reset),
    .value (_col_1_n_w3_add_w5_value)
  );
  W6 col_1_n_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1062:64
    .clock (clock),
    .reset (reset),
    .value (_col_1_n_w6_value)
  );
  W2_sub_W6 col_1_n_w2_sub_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1063:85
    .clock (clock),
    .reset (reset),
    .value (_col_1_n_w2_sub_w6_value)
  );
  W2_add_W6 col_1_n_w2_add_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1064:85
    .clock (clock),
    .reset (reset),
    .value (_col_1_n_w2_add_w6_value)
  );
  SHL_8 col_1_n_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1065:83
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_shr_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:623:87
    .z     (_col_1_n_x1_0_z)
  );
  SHL_8 col_1_n_t0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1066:83
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_shr_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:231:87
    .z     (_col_1_n_t0_0_z)
  );
  ADD col_1_n_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1067:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_t0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1066:83
    .y     (_col_1_n_c8192_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1055:73
    .z     (_col_1_n_x0_0_z)
  );
  dup_2 col_1_d_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1068:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1067:100
    .y     (_col_1_d_x0_0_y),
    .z     (_col_1_d_x0_0_z)
  );
  dup_2 col_1_d_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1069:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1065:83
    .y     (_col_1_d_x1_0_y),
    .z     (_col_1_d_x1_0_z)
  );
  dup_2 col_1_d_x2_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1070:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_shr_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:819:87
    .y     (_col_1_d_x2_0_y),
    .z     (_col_1_d_x2_0_z)
  );
  dup_2 col_1_d_x3_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1071:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_shr_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:427:87
    .y     (_col_1_d_x3_0_y),
    .z     (_col_1_d_x3_0_z)
  );
  dup_2 col_1_d_x4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1072:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_shr_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:329:87
    .y     (_col_1_d_x4_0_y),
    .z     (_col_1_d_x4_0_z)
  );
  dup_2 col_1_d_x5_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1073:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_shr_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:917:87
    .y     (_col_1_d_x5_0_y),
    .z     (_col_1_d_x5_0_z)
  );
  dup_2 col_1_d_x6_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1074:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_shr_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:721:87
    .y     (_col_1_d_x6_0_y),
    .z     (_col_1_d_x6_0_z)
  );
  dup_2 col_1_d_x7_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1075:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_shr_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:525:87
    .y     (_col_1_d_x7_0_y),
    .z     (_col_1_d_x7_0_z)
  );
  ADD col_1_n_u8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1076:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_129_1988_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2006:118
    .y     (_col_1_d_x5_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1073:100
    .z     (_col_1_n_u8_0_z)
  );
  MUL col_1_n_v8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1077:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1056:64
    .y     (_col_1_n_u8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1076:100
    .z     (_col_1_n_v8_0_z)
  );
  ADD col_1_n_x8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1078:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_v8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1077:100
    .y     (_col_1_n_c4_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1048:70
    .z     (_col_1_n_x8_0_z)
  );
  dup_2 col_1_d_x8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1079:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1078:100
    .y     (_col_1_d_x8_0_y),
    .z     (_col_1_d_x8_0_z)
  );
  MUL col_1_n_u4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1080:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_w1_sub_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1057:85
    .y     (_col_1_d_x4_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1072:100
    .z     (_col_1_n_u4_1_z)
  );
  ADD col_1_n_v4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1081:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x8_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1079:100
    .y     (_delay_INT16_262_1987_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2005:118
    .z     (_col_1_n_v4_1_z)
  );
  SHR_3 col_1_n_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1082:83
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_v4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1081:100
    .z     (_col_1_n_x4_1_z)
  );
  dup_2 col_1_d_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1083:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1082:83
    .y     (_col_1_d_x4_1_y),
    .z     (_col_1_d_x4_1_z)
  );
  MUL col_1_n_u5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1084:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_w1_add_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1058:85
    .y     (_col_1_d_x5_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1073:100
    .z     (_col_1_n_u5_1_z)
  );
  SUB col_1_n_v5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1085:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1079:100
    .y     (_delay_INT16_90_1986_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2004:114
    .z     (_col_1_n_v5_1_z)
  );
  SHR_3 col_1_n_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1086:83
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_v5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1085:100
    .z     (_col_1_n_x5_1_z)
  );
  dup_2 col_1_d_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1087:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1086:83
    .y     (_col_1_d_x5_1_y),
    .z     (_col_1_d_x5_1_z)
  );
  ADD col_1_n_u8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1088:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_88_1985_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2003:114
    .y     (_col_1_d_x7_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1075:100
    .z     (_col_1_n_u8_1_z)
  );
  MUL col_1_n_v8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1089:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_w3_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1059:64
    .y     (_col_1_n_u8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1088:100
    .z     (_col_1_n_v8_1_z)
  );
  ADD col_1_n_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1090:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_v8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1089:100
    .y     (_col_1_n_c4_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1049:70
    .z     (_col_1_n_x8_1_z)
  );
  dup_2 col_1_d_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1091:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1090:100
    .y     (_col_1_d_x8_1_y),
    .z     (_col_1_d_x8_1_z)
  );
  MUL col_1_n_u6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1092:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_w3_sub_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1060:85
    .y     (_col_1_d_x6_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1074:100
    .z     (_col_1_n_u6_1_z)
  );
  SUB col_1_n_v6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1093:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x8_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1091:100
    .y     (_delay_INT16_191_1983_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2001:118
    .z     (_col_1_n_v6_1_z)
  );
  SHR_3 col_1_n_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1094:83
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_v6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1093:100
    .z     (_col_1_n_x6_1_z)
  );
  dup_2 col_1_d_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1095:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1094:83
    .y     (_col_1_d_x6_1_y),
    .z     (_col_1_d_x6_1_z)
  );
  MUL col_1_n_u7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1096:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_w3_add_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1061:85
    .y     (_col_1_d_x7_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1075:100
    .z     (_col_1_n_u7_1_z)
  );
  SUB col_1_n_v7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1097:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1091:100
    .y     (_delay_INT16_102_1982_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2000:118
    .z     (_col_1_n_v7_1_z)
  );
  SHR_3 col_1_n_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1098:83
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_v7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1097:100
    .z     (_col_1_n_x7_1_z)
  );
  dup_2 col_1_d_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1099:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1098:83
    .y     (_col_1_d_x7_1_y),
    .z     (_col_1_d_x7_1_z)
  );
  ADD col_1_n_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1100:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x0_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1068:100
    .y     (_delay_INT16_131_1981_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1999:118
    .z     (_col_1_n_x8_2_z)
  );
  dup_2 col_1_d_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1101:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1100:100
    .y     (_col_1_d_x8_2_y),
    .z     (_col_1_d_x8_2_z)
  );
  SUB col_1_n_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1102:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1068:100
    .y     (_delay_INT16_131_1979_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1997:118
    .z     (_col_1_n_x0_1_z)
  );
  dup_2 col_1_d_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1103:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1102:100
    .y     (_col_1_d_x0_1_y),
    .z     (_col_1_d_x0_1_z)
  );
  ADD col_1_n_u1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1104:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_62_2052_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2070:114
    .y     (_col_1_d_x2_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1070:100
    .z     (_col_1_n_u1_1_z)
  );
  MUL col_1_n_v1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1105:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1062:64
    .y     (_col_1_n_u1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1104:100
    .z     (_col_1_n_v1_1_z)
  );
  ADD col_1_n_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1106:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_v1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1105:100
    .y     (_col_1_n_c4_2_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1050:70
    .z     (_col_1_n_x1_1_z)
  );
  dup_2 col_1_d_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1107:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1106:100
    .y     (_col_1_d_x1_1_y),
    .z     (_col_1_d_x1_1_z)
  );
  MUL col_1_n_u2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1108:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_w2_add_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1064:85
    .y     (_col_1_d_x2_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1070:100
    .z     (_col_1_n_u2_1_z)
  );
  SUB col_1_n_v2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1109:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x1_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1107:100
    .y     (_delay_INT16_109_1977_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1995:118
    .z     (_col_1_n_v2_1_z)
  );
  SHR_3 col_1_n_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1110:83
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_v2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1109:100
    .z     (_col_1_n_x2_1_z)
  );
  dup_2 col_1_d_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1111:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1110:83
    .y     (_col_1_d_x2_1_y),
    .z     (_col_1_d_x2_1_z)
  );
  MUL col_1_n_u3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1112:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_w2_sub_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1063:85
    .y     (_col_1_d_x3_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1071:100
    .z     (_col_1_n_u3_1_z)
  );
  ADD col_1_n_v3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1113:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1107:100
    .y     (_delay_INT16_259_1984_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2002:118
    .z     (_col_1_n_v3_1_z)
  );
  SHR_3 col_1_n_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1114:83
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_v3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1113:100
    .z     (_col_1_n_x3_1_z)
  );
  dup_2 col_1_d_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1115:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1114:83
    .y     (_col_1_d_x3_1_y),
    .z     (_col_1_d_x3_1_z)
  );
  ADD col_1_n_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1116:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x4_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1083:100
    .y     (_delay_INT16_64_2020_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2038:114
    .z     (_col_1_n_x1_2_z)
  );
  dup_2 col_1_d_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1117:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1116:100
    .y     (_col_1_d_x1_2_y),
    .z     (_col_1_d_x1_2_z)
  );
  SUB col_1_n_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1118:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1083:100
    .y     (_delay_INT16_64_1976_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1994:114
    .z     (_col_1_n_x4_2_z)
  );
  dup_2 col_1_d_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1119:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1118:100
    .y     (_col_1_d_x4_2_y),
    .z     (_col_1_d_x4_2_z)
  );
  ADD col_1_n_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1120:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x5_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1087:100
    .y     (_delay_INT16_10_1975_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1993:114
    .z     (_col_1_n_x6_2_z)
  );
  dup_2 col_1_d_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1121:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1120:100
    .y     (_col_1_d_x6_2_y),
    .z     (_col_1_d_x6_2_z)
  );
  SUB col_1_n_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1122:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1087:100
    .y     (_delay_INT16_10_1974_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1992:114
    .z     (_col_1_n_x5_2_z)
  );
  dup_2 col_1_d_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1123:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1122:100
    .y     (_col_1_d_x5_2_y),
    .z     (_col_1_d_x5_2_z)
  );
  ADD col_1_n_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1124:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x8_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1101:100
    .y     (_delay_INT16_27_1973_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1991:114
    .z     (_col_1_n_x7_2_z)
  );
  dup_2 col_1_d_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1125:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1124:100
    .y     (_col_1_d_x7_2_y),
    .z     (_col_1_d_x7_2_z)
  );
  SUB col_1_n_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1126:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1101:100
    .y     (_delay_INT16_27_1972_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1990:114
    .z     (_col_1_n_x8_3_z)
  );
  dup_2 col_1_d_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1127:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1126:100
    .y     (_col_1_d_x8_3_y),
    .z     (_col_1_d_x8_3_z)
  );
  ADD col_1_n_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1128:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_45_1970_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1988:114
    .y     (_col_1_d_x2_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1111:100
    .z     (_col_1_n_x3_2_z)
  );
  dup_2 col_1_d_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1129:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1128:100
    .y     (_col_1_d_x3_2_y),
    .z     (_col_1_d_x3_2_z)
  );
  SUB col_1_n_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1130:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_45_1969_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1987:114
    .y     (_col_1_d_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1111:100
    .z     (_col_1_n_x0_2_z)
  );
  dup_2 col_1_d_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1131:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1130:100
    .y     (_col_1_d_x0_2_y),
    .z     (_col_1_d_x0_2_z)
  );
  ADD col_1_n_u2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1132:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_2_1968_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1986:110
    .y     (_col_1_d_x5_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1123:100
    .z     (_col_1_n_u2_2_z)
  );
  MUL col_1_n_v2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1133:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_c181_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1053:76
    .y     (_col_1_n_u2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1132:100
    .z     (_col_1_n_v2_2_z)
  );
  ADD col_1_n_w2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1134:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_v2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1133:100
    .y     (_col_1_n_c128_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1051:76
    .z     (_col_1_n_w2_2_z)
  );
  SHR_8 col_1_n_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1135:83
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_w2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1134:100
    .z     (_col_1_n_x2_2_z)
  );
  dup_2 col_1_d_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1136:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1135:83
    .y     (_col_1_d_x2_2_y),
    .z     (_col_1_d_x2_2_z)
  );
  SUB col_1_n_u4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1137:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_2_2081_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2099:110
    .y     (_col_1_d_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1123:100
    .z     (_col_1_n_u4_3_z)
  );
  MUL col_1_n_v4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1138:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_c181_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1054:76
    .y     (_col_1_n_u4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1137:100
    .z     (_col_1_n_v4_3_z)
  );
  ADD col_1_n_w4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1139:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_v4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1138:100
    .y     (_col_1_n_c128_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1052:76
    .z     (_col_1_n_w4_3_z)
  );
  SHR_8 col_1_n_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1140:83
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_w4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1139:100
    .z     (_col_1_n_x4_3_z)
  );
  dup_2 col_1_d_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1141:100
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1140:83
    .y     (_col_1_d_x4_3_y),
    .z     (_col_1_d_x4_3_z)
  );
  ADD col_1_n_tmp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1142:105
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x7_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1125:100
    .y     (_delay_INT16_1_1966_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1984:110
    .z     (_col_1_n_tmp_0_z)
  );
  SHR_14 col_1_n_val_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1143:87
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_tmp_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1142:105
    .z     (_col_1_n_val_0_z)
  );
  CLIP col_1_n_clp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1144:87
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_val_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1143:87
    .z     (n_out_0_1_x)
  );
  ADD col_1_n_tmp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1145:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_190_1965_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1983:118
    .y     (_col_1_d_x2_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1136:100
    .z     (_col_1_n_tmp_1_z)
  );
  SHR_14 col_1_n_val_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1146:87
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_tmp_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1145:105
    .z     (_col_1_n_val_1_z)
  );
  CLIP col_1_n_clp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1147:87
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_val_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1146:87
    .z     (n_out_1_1_x)
  );
  ADD col_1_n_tmp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1148:105
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x0_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1131:100
    .y     (_delay_INT16_19_2324_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2342:114
    .z     (_col_1_n_tmp_2_z)
  );
  SHR_14 col_1_n_val_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1149:87
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_tmp_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1148:105
    .z     (_col_1_n_val_2_z)
  );
  CLIP col_1_n_clp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1150:87
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_val_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1149:87
    .z     (n_out_2_1_x)
  );
  ADD col_1_n_tmp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1151:105
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x8_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1127:100
    .y     (_delay_INT16_73_1964_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1982:114
    .z     (_col_1_n_tmp_3_z)
  );
  SHR_14 col_1_n_val_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1152:87
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_tmp_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1151:105
    .z     (_col_1_n_val_3_z)
  );
  CLIP col_1_n_clp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1153:87
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_val_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1152:87
    .z     (n_out_3_1_x)
  );
  SUB col_1_n_tmp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1154:105
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1127:100
    .y     (_delay_INT16_73_2111_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2129:114
    .z     (_col_1_n_tmp_4_z)
  );
  SHR_14 col_1_n_val_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1155:87
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_tmp_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1154:105
    .z     (_col_1_n_val_4_z)
  );
  CLIP col_1_n_clp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1156:87
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_val_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1155:87
    .z     (n_out_4_1_x)
  );
  SUB col_1_n_tmp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1157:105
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1131:100
    .y     (_delay_INT16_19_1963_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1981:114
    .z     (_col_1_n_tmp_5_z)
  );
  SHR_14 col_1_n_val_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1158:87
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_tmp_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1157:105
    .z     (_col_1_n_val_5_z)
  );
  CLIP col_1_n_clp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1159:87
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_val_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1158:87
    .z     (n_out_5_1_x)
  );
  SUB col_1_n_tmp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1160:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_190_1962_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1980:118
    .y     (_col_1_d_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1136:100
    .z     (_col_1_n_tmp_6_z)
  );
  SHR_14 col_1_n_val_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1161:87
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_tmp_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1160:105
    .z     (_col_1_n_val_6_z)
  );
  CLIP col_1_n_clp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1162:87
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_val_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1161:87
    .z     (n_out_6_1_x)
  );
  SUB col_1_n_tmp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1163:105
    .clock (clock),
    .reset (reset),
    .x     (_col_1_d_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1125:100
    .y     (_delay_INT16_1_1961_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1979:110
    .z     (_col_1_n_tmp_7_z)
  );
  SHR_14 col_1_n_val_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1164:87
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_tmp_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1163:105
    .z     (_col_1_n_val_7_z)
  );
  CLIP col_1_n_clp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1165:87
    .clock (clock),
    .reset (reset),
    .x     (_col_1_n_val_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1164:87
    .z     (n_out_7_1_x)
  );
  C4 col_2_n_c4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1166:70
    .clock (clock),
    .reset (reset),
    .value (_col_2_n_c4_0_value)
  );
  C4 col_2_n_c4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1167:70
    .clock (clock),
    .reset (reset),
    .value (_col_2_n_c4_1_value)
  );
  C4 col_2_n_c4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1168:70
    .clock (clock),
    .reset (reset),
    .value (_col_2_n_c4_2_value)
  );
  C128 col_2_n_c128_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1169:76
    .clock (clock),
    .reset (reset),
    .value (_col_2_n_c128_0_value)
  );
  C128 col_2_n_c128_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1170:76
    .clock (clock),
    .reset (reset),
    .value (_col_2_n_c128_1_value)
  );
  C181 col_2_n_c181_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1171:76
    .clock (clock),
    .reset (reset),
    .value (_col_2_n_c181_0_value)
  );
  C181 col_2_n_c181_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1172:76
    .clock (clock),
    .reset (reset),
    .value (_col_2_n_c181_1_value)
  );
  C8192 col_2_n_c8192 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1173:73
    .clock (clock),
    .reset (reset),
    .value (_col_2_n_c8192_value)
  );
  W7 col_2_n_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1174:64
    .clock (clock),
    .reset (reset),
    .value (_col_2_n_w7_value)
  );
  W1_sub_W7 col_2_n_w1_sub_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1175:85
    .clock (clock),
    .reset (reset),
    .value (_col_2_n_w1_sub_w7_value)
  );
  W1_add_W7 col_2_n_w1_add_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1176:85
    .clock (clock),
    .reset (reset),
    .value (_col_2_n_w1_add_w7_value)
  );
  W3 col_2_n_w3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1177:64
    .clock (clock),
    .reset (reset),
    .value (_col_2_n_w3_value)
  );
  W3_sub_W5 col_2_n_w3_sub_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1178:85
    .clock (clock),
    .reset (reset),
    .value (_col_2_n_w3_sub_w5_value)
  );
  W3_add_W5 col_2_n_w3_add_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1179:85
    .clock (clock),
    .reset (reset),
    .value (_col_2_n_w3_add_w5_value)
  );
  W6 col_2_n_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1180:64
    .clock (clock),
    .reset (reset),
    .value (_col_2_n_w6_value)
  );
  W2_sub_W6 col_2_n_w2_sub_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1181:85
    .clock (clock),
    .reset (reset),
    .value (_col_2_n_w2_sub_w6_value)
  );
  W2_add_W6 col_2_n_w2_add_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1182:85
    .clock (clock),
    .reset (reset),
    .value (_col_2_n_w2_add_w6_value)
  );
  SHL_8 col_2_n_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1183:83
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_shr_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:625:87
    .z     (_col_2_n_x1_0_z)
  );
  SHL_8 col_2_n_t0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1184:83
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_shr_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:233:87
    .z     (_col_2_n_t0_0_z)
  );
  ADD col_2_n_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1185:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_t0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1184:83
    .y     (_col_2_n_c8192_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1173:73
    .z     (_col_2_n_x0_0_z)
  );
  dup_2 col_2_d_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1186:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1185:100
    .y     (_col_2_d_x0_0_y),
    .z     (_col_2_d_x0_0_z)
  );
  dup_2 col_2_d_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1187:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1183:83
    .y     (_col_2_d_x1_0_y),
    .z     (_col_2_d_x1_0_z)
  );
  dup_2 col_2_d_x2_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1188:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_shr_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:821:87
    .y     (_col_2_d_x2_0_y),
    .z     (_col_2_d_x2_0_z)
  );
  dup_2 col_2_d_x3_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1189:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_shr_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:429:87
    .y     (_col_2_d_x3_0_y),
    .z     (_col_2_d_x3_0_z)
  );
  dup_2 col_2_d_x4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1190:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_shr_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:331:87
    .y     (_col_2_d_x4_0_y),
    .z     (_col_2_d_x4_0_z)
  );
  dup_2 col_2_d_x5_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1191:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_shr_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:919:87
    .y     (_col_2_d_x5_0_y),
    .z     (_col_2_d_x5_0_z)
  );
  dup_2 col_2_d_x6_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1192:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_shr_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:723:87
    .y     (_col_2_d_x6_0_y),
    .z     (_col_2_d_x6_0_z)
  );
  dup_2 col_2_d_x7_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1193:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_shr_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:527:87
    .y     (_col_2_d_x7_0_y),
    .z     (_col_2_d_x7_0_z)
  );
  ADD col_2_n_u8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1194:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_34_1959_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1977:114
    .y     (_col_2_d_x5_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1191:100
    .z     (_col_2_n_u8_0_z)
  );
  MUL col_2_n_v8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1195:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1174:64
    .y     (_col_2_n_u8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1194:100
    .z     (_col_2_n_v8_0_z)
  );
  ADD col_2_n_x8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1196:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_v8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1195:100
    .y     (_col_2_n_c4_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1166:70
    .z     (_col_2_n_x8_0_z)
  );
  dup_2 col_2_d_x8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1197:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1196:100
    .y     (_col_2_d_x8_0_y),
    .z     (_col_2_d_x8_0_z)
  );
  MUL col_2_n_u4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1198:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_w1_sub_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1175:85
    .y     (_col_2_d_x4_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1190:100
    .z     (_col_2_n_u4_1_z)
  );
  ADD col_2_n_v4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1199:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_d_x8_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1197:100
    .y     (_delay_INT16_112_1958_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1976:118
    .z     (_col_2_n_v4_1_z)
  );
  SHR_3 col_2_n_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1200:83
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_v4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1199:100
    .z     (_col_2_n_x4_1_z)
  );
  dup_2 col_2_d_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1201:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1200:83
    .y     (_col_2_d_x4_1_y),
    .z     (_col_2_d_x4_1_z)
  );
  MUL col_2_n_u5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1202:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_w1_add_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1176:85
    .y     (_col_2_d_x5_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1191:100
    .z     (_col_2_n_u5_1_z)
  );
  SUB col_2_n_v5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1203:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_d_x8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1197:100
    .y     (_delay_INT16_68_1957_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1975:114
    .z     (_col_2_n_v5_1_z)
  );
  SHR_3 col_2_n_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1204:83
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_v5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1203:100
    .z     (_col_2_n_x5_1_z)
  );
  dup_2 col_2_d_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1205:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1204:83
    .y     (_col_2_d_x5_1_y),
    .z     (_col_2_d_x5_1_z)
  );
  ADD col_2_n_u8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1206:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_1_2294_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2312:110
    .y     (_col_2_d_x7_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1193:100
    .z     (_col_2_n_u8_1_z)
  );
  MUL col_2_n_v8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1207:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_w3_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1177:64
    .y     (_col_2_n_u8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1206:100
    .z     (_col_2_n_v8_1_z)
  );
  ADD col_2_n_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1208:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_v8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1207:100
    .y     (_col_2_n_c4_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1167:70
    .z     (_col_2_n_x8_1_z)
  );
  dup_2 col_2_d_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1209:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1208:100
    .y     (_col_2_d_x8_1_y),
    .z     (_col_2_d_x8_1_z)
  );
  MUL col_2_n_u6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1210:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_w3_sub_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1178:85
    .y     (_col_2_d_x6_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1192:100
    .z     (_col_2_n_u6_1_z)
  );
  SUB col_2_n_v6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1211:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_d_x8_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1209:100
    .y     (_delay_INT16_50_2056_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2074:114
    .z     (_col_2_n_v6_1_z)
  );
  SHR_3 col_2_n_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1212:83
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_v6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1211:100
    .z     (_col_2_n_x6_1_z)
  );
  dup_2 col_2_d_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1213:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1212:83
    .y     (_col_2_d_x6_1_y),
    .z     (_col_2_d_x6_1_z)
  );
  MUL col_2_n_u7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1214:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_w3_add_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1179:85
    .y     (_col_2_d_x7_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1193:100
    .z     (_col_2_n_u7_1_z)
  );
  SUB col_2_n_v7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1215:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_d_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1209:100
    .y     (_delay_INT16_131_1956_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1974:118
    .z     (_col_2_n_v7_1_z)
  );
  SHR_3 col_2_n_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1216:83
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_v7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1215:100
    .z     (_col_2_n_x7_1_z)
  );
  dup_2 col_2_d_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1217:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1216:83
    .y     (_col_2_d_x7_1_y),
    .z     (_col_2_d_x7_1_z)
  );
  ADD col_2_n_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1218:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_213_1955_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1973:118
    .y     (_col_2_d_x1_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1187:100
    .z     (_col_2_n_x8_2_z)
  );
  dup_2 col_2_d_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1219:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1218:100
    .y     (_col_2_d_x8_2_y),
    .z     (_col_2_d_x8_2_z)
  );
  SUB col_2_n_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1220:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_213_1989_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2007:118
    .y     (_col_2_d_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1187:100
    .z     (_col_2_n_x0_1_z)
  );
  dup_2 col_2_d_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1221:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1220:100
    .y     (_col_2_d_x0_1_y),
    .z     (_col_2_d_x0_1_z)
  );
  ADD col_2_n_u1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1222:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_66_1954_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1972:114
    .y     (_col_2_d_x2_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1188:100
    .z     (_col_2_n_u1_1_z)
  );
  MUL col_2_n_v1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1223:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1180:64
    .y     (_col_2_n_u1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1222:100
    .z     (_col_2_n_v1_1_z)
  );
  ADD col_2_n_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1224:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_v1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1223:100
    .y     (_col_2_n_c4_2_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1168:70
    .z     (_col_2_n_x1_1_z)
  );
  dup_2 col_2_d_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1225:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1224:100
    .y     (_col_2_d_x1_1_y),
    .z     (_col_2_d_x1_1_z)
  );
  MUL col_2_n_u2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1226:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_w2_add_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1182:85
    .y     (_col_2_d_x2_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1188:100
    .z     (_col_2_n_u2_1_z)
  );
  SUB col_2_n_v2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1227:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_d_x1_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1225:100
    .y     (_delay_INT16_156_2021_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2039:118
    .z     (_col_2_n_v2_1_z)
  );
  SHR_3 col_2_n_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1228:83
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_v2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1227:100
    .z     (_col_2_n_x2_1_z)
  );
  dup_2 col_2_d_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1229:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1228:83
    .y     (_col_2_d_x2_1_y),
    .z     (_col_2_d_x2_1_z)
  );
  MUL col_2_n_u3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1230:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_w2_sub_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1181:85
    .y     (_col_2_d_x3_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1189:100
    .z     (_col_2_n_u3_1_z)
  );
  ADD col_2_n_v3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1231:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_d_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1225:100
    .y     (_delay_INT16_168_1953_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1971:118
    .z     (_col_2_n_v3_1_z)
  );
  SHR_3 col_2_n_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1232:83
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_v3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1231:100
    .z     (_col_2_n_x3_1_z)
  );
  dup_2 col_2_d_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1233:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1232:83
    .y     (_col_2_d_x3_1_y),
    .z     (_col_2_d_x3_1_z)
  );
  ADD col_2_n_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1234:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_78_2205_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2223:114
    .y     (_col_2_d_x6_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1213:100
    .z     (_col_2_n_x1_2_z)
  );
  dup_2 col_2_d_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1235:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1234:100
    .y     (_col_2_d_x1_2_y),
    .z     (_col_2_d_x1_2_z)
  );
  SUB col_2_n_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1236:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_78_2091_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2109:114
    .y     (_col_2_d_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1213:100
    .z     (_col_2_n_x4_2_z)
  );
  dup_2 col_2_d_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1237:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1236:100
    .y     (_col_2_d_x4_2_y),
    .z     (_col_2_d_x4_2_z)
  );
  ADD col_2_n_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1238:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_64_2231_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2249:114
    .y     (_col_2_d_x7_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1217:100
    .z     (_col_2_n_x6_2_z)
  );
  dup_2 col_2_d_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1239:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1238:100
    .y     (_col_2_d_x6_2_y),
    .z     (_col_2_d_x6_2_z)
  );
  SUB col_2_n_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1240:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_64_1952_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1970:114
    .y     (_col_2_d_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1217:100
    .z     (_col_2_n_x5_2_z)
  );
  dup_2 col_2_d_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1241:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1240:100
    .y     (_col_2_d_x5_2_y),
    .z     (_col_2_d_x5_2_z)
  );
  ADD col_2_n_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1242:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_d_x8_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1219:100
    .y     (_delay_INT16_75_2268_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2286:114
    .z     (_col_2_n_x7_2_z)
  );
  dup_2 col_2_d_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1243:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1242:100
    .y     (_col_2_d_x7_2_y),
    .z     (_col_2_d_x7_2_z)
  );
  SUB col_2_n_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1244:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_d_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1219:100
    .y     (_delay_INT16_75_1951_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1969:114
    .z     (_col_2_n_x8_3_z)
  );
  dup_2 col_2_d_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1245:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1244:100
    .y     (_col_2_d_x8_3_y),
    .z     (_col_2_d_x8_3_z)
  );
  ADD col_2_n_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1246:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_66_1950_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1968:114
    .y     (_col_2_d_x2_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1229:100
    .z     (_col_2_n_x3_2_z)
  );
  dup_2 col_2_d_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1247:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1246:100
    .y     (_col_2_d_x3_2_y),
    .z     (_col_2_d_x3_2_z)
  );
  SUB col_2_n_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1248:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_66_2121_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2139:114
    .y     (_col_2_d_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1229:100
    .z     (_col_2_n_x0_2_z)
  );
  dup_2 col_2_d_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1249:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1248:100
    .y     (_col_2_d_x0_2_y),
    .z     (_col_2_d_x0_2_z)
  );
  ADD col_2_n_u2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1250:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_d_x4_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1237:100
    .y     (_delay_INT16_90_2010_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2028:114
    .z     (_col_2_n_u2_2_z)
  );
  MUL col_2_n_v2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1251:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_c181_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1171:76
    .y     (_col_2_n_u2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1250:100
    .z     (_col_2_n_v2_2_z)
  );
  ADD col_2_n_w2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1252:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_v2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1251:100
    .y     (_col_2_n_c128_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1169:76
    .z     (_col_2_n_w2_2_z)
  );
  SHR_8 col_2_n_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1253:83
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_w2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1252:100
    .z     (_col_2_n_x2_2_z)
  );
  dup_2 col_2_d_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1254:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1253:83
    .y     (_col_2_d_x2_2_y),
    .z     (_col_2_d_x2_2_z)
  );
  SUB col_2_n_u4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1255:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_d_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1237:100
    .y     (_delay_INT16_90_1946_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1964:114
    .z     (_col_2_n_u4_3_z)
  );
  MUL col_2_n_v4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1256:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_c181_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1172:76
    .y     (_col_2_n_u4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1255:100
    .z     (_col_2_n_v4_3_z)
  );
  ADD col_2_n_w4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1257:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_v4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1256:100
    .y     (_col_2_n_c128_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1170:76
    .z     (_col_2_n_w4_3_z)
  );
  SHR_8 col_2_n_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1258:83
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_w4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1257:100
    .z     (_col_2_n_x4_3_z)
  );
  dup_2 col_2_d_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1259:100
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1258:83
    .y     (_col_2_d_x4_3_y),
    .z     (_col_2_d_x4_3_z)
  );
  ADD col_2_n_tmp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1260:105
    .clock (clock),
    .reset (reset),
    .x     (_col_2_d_x7_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1243:100
    .y     (_delay_INT16_122_1945_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1963:118
    .z     (_col_2_n_tmp_0_z)
  );
  SHR_14 col_2_n_val_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1261:87
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_tmp_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1260:105
    .z     (_col_2_n_val_0_z)
  );
  CLIP col_2_n_clp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1262:87
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_val_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1261:87
    .z     (n_out_0_2_x)
  );
  ADD col_2_n_tmp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1263:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_121_1944_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1962:118
    .y     (_col_2_d_x2_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1254:100
    .z     (_col_2_n_tmp_1_z)
  );
  SHR_14 col_2_n_val_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1264:87
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_tmp_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1263:105
    .z     (_col_2_n_val_1_z)
  );
  CLIP col_2_n_clp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1265:87
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_val_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1264:87
    .z     (n_out_1_2_x)
  );
  ADD col_2_n_tmp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1266:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_110_1943_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1961:118
    .y     (_col_2_d_x4_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1259:100
    .z     (_col_2_n_tmp_2_z)
  );
  SHR_14 col_2_n_val_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1267:87
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_tmp_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1266:105
    .z     (_col_2_n_val_2_z)
  );
  CLIP col_2_n_clp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1268:87
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_val_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1267:87
    .z     (n_out_2_2_x)
  );
  ADD col_2_n_tmp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1269:105
    .clock (clock),
    .reset (reset),
    .x     (_col_2_d_x8_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1245:100
    .y     (_delay_INT16_145_1942_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1960:118
    .z     (_col_2_n_tmp_3_z)
  );
  SHR_14 col_2_n_val_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1270:87
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_tmp_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1269:105
    .z     (_col_2_n_val_3_z)
  );
  CLIP col_2_n_clp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1271:87
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_val_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1270:87
    .z     (n_out_3_2_x)
  );
  SUB col_2_n_tmp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1272:105
    .clock (clock),
    .reset (reset),
    .x     (_col_2_d_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1245:100
    .y     (_delay_INT16_145_2015_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2033:118
    .z     (_col_2_n_tmp_4_z)
  );
  SHR_14 col_2_n_val_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1273:87
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_tmp_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1272:105
    .z     (_col_2_n_val_4_z)
  );
  CLIP col_2_n_clp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1274:87
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_val_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1273:87
    .z     (n_out_4_2_x)
  );
  SUB col_2_n_tmp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1275:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_110_1941_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1959:118
    .y     (_col_2_d_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1259:100
    .z     (_col_2_n_tmp_5_z)
  );
  SHR_14 col_2_n_val_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1276:87
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_tmp_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1275:105
    .z     (_col_2_n_val_5_z)
  );
  CLIP col_2_n_clp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1277:87
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_val_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1276:87
    .z     (n_out_5_2_x)
  );
  SUB col_2_n_tmp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1278:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_121_1940_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1958:118
    .y     (_col_2_d_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1254:100
    .z     (_col_2_n_tmp_6_z)
  );
  SHR_14 col_2_n_val_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1279:87
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_tmp_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1278:105
    .z     (_col_2_n_val_6_z)
  );
  CLIP col_2_n_clp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1280:87
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_val_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1279:87
    .z     (n_out_6_2_x)
  );
  SUB col_2_n_tmp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1281:105
    .clock (clock),
    .reset (reset),
    .x     (_col_2_d_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1243:100
    .y     (_delay_INT16_122_1939_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1957:118
    .z     (_col_2_n_tmp_7_z)
  );
  SHR_14 col_2_n_val_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1282:87
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_tmp_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1281:105
    .z     (_col_2_n_val_7_z)
  );
  CLIP col_2_n_clp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1283:87
    .clock (clock),
    .reset (reset),
    .x     (_col_2_n_val_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1282:87
    .z     (n_out_7_2_x)
  );
  C4 col_3_n_c4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1284:70
    .clock (clock),
    .reset (reset),
    .value (_col_3_n_c4_0_value)
  );
  C4 col_3_n_c4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1285:70
    .clock (clock),
    .reset (reset),
    .value (_col_3_n_c4_1_value)
  );
  C4 col_3_n_c4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1286:70
    .clock (clock),
    .reset (reset),
    .value (_col_3_n_c4_2_value)
  );
  C128 col_3_n_c128_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1287:76
    .clock (clock),
    .reset (reset),
    .value (_col_3_n_c128_0_value)
  );
  C128 col_3_n_c128_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1288:76
    .clock (clock),
    .reset (reset),
    .value (_col_3_n_c128_1_value)
  );
  C181 col_3_n_c181_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1289:76
    .clock (clock),
    .reset (reset),
    .value (_col_3_n_c181_0_value)
  );
  C181 col_3_n_c181_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1290:76
    .clock (clock),
    .reset (reset),
    .value (_col_3_n_c181_1_value)
  );
  C8192 col_3_n_c8192 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1291:73
    .clock (clock),
    .reset (reset),
    .value (_col_3_n_c8192_value)
  );
  W7 col_3_n_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1292:64
    .clock (clock),
    .reset (reset),
    .value (_col_3_n_w7_value)
  );
  W1_sub_W7 col_3_n_w1_sub_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1293:85
    .clock (clock),
    .reset (reset),
    .value (_col_3_n_w1_sub_w7_value)
  );
  W1_add_W7 col_3_n_w1_add_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1294:85
    .clock (clock),
    .reset (reset),
    .value (_col_3_n_w1_add_w7_value)
  );
  W3 col_3_n_w3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1295:64
    .clock (clock),
    .reset (reset),
    .value (_col_3_n_w3_value)
  );
  W3_sub_W5 col_3_n_w3_sub_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1296:85
    .clock (clock),
    .reset (reset),
    .value (_col_3_n_w3_sub_w5_value)
  );
  W3_add_W5 col_3_n_w3_add_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1297:85
    .clock (clock),
    .reset (reset),
    .value (_col_3_n_w3_add_w5_value)
  );
  W6 col_3_n_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1298:64
    .clock (clock),
    .reset (reset),
    .value (_col_3_n_w6_value)
  );
  W2_sub_W6 col_3_n_w2_sub_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1299:85
    .clock (clock),
    .reset (reset),
    .value (_col_3_n_w2_sub_w6_value)
  );
  W2_add_W6 col_3_n_w2_add_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1300:85
    .clock (clock),
    .reset (reset),
    .value (_col_3_n_w2_add_w6_value)
  );
  SHL_8 col_3_n_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1301:83
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_shr_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:627:87
    .z     (_col_3_n_x1_0_z)
  );
  SHL_8 col_3_n_t0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1302:83
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_shr_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:235:87
    .z     (_col_3_n_t0_0_z)
  );
  ADD col_3_n_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1303:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_t0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1302:83
    .y     (_col_3_n_c8192_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1291:73
    .z     (_col_3_n_x0_0_z)
  );
  dup_2 col_3_d_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1304:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1303:100
    .y     (_col_3_d_x0_0_y),
    .z     (_col_3_d_x0_0_z)
  );
  dup_2 col_3_d_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1305:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1301:83
    .y     (_col_3_d_x1_0_y),
    .z     (_col_3_d_x1_0_z)
  );
  dup_2 col_3_d_x2_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1306:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_shr_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:823:87
    .y     (_col_3_d_x2_0_y),
    .z     (_col_3_d_x2_0_z)
  );
  dup_2 col_3_d_x3_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1307:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_shr_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:431:87
    .y     (_col_3_d_x3_0_y),
    .z     (_col_3_d_x3_0_z)
  );
  dup_2 col_3_d_x4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1308:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_shr_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:333:87
    .y     (_col_3_d_x4_0_y),
    .z     (_col_3_d_x4_0_z)
  );
  dup_2 col_3_d_x5_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1309:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_shr_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:921:87
    .y     (_col_3_d_x5_0_y),
    .z     (_col_3_d_x5_0_z)
  );
  dup_2 col_3_d_x6_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1310:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_shr_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:725:87
    .y     (_col_3_d_x6_0_y),
    .z     (_col_3_d_x6_0_z)
  );
  dup_2 col_3_d_x7_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1311:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_shr_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:529:87
    .y     (_col_3_d_x7_0_y),
    .z     (_col_3_d_x7_0_z)
  );
  ADD col_3_n_u8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1312:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_65_1937_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1955:114
    .y     (_col_3_d_x5_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1309:100
    .z     (_col_3_n_u8_0_z)
  );
  MUL col_3_n_v8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1313:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1292:64
    .y     (_col_3_n_u8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1312:100
    .z     (_col_3_n_v8_0_z)
  );
  ADD col_3_n_x8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1314:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_v8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1313:100
    .y     (_col_3_n_c4_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1284:70
    .z     (_col_3_n_x8_0_z)
  );
  dup_2 col_3_d_x8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1315:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1314:100
    .y     (_col_3_d_x8_0_y),
    .z     (_col_3_d_x8_0_z)
  );
  MUL col_3_n_u4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1316:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_w1_sub_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1293:85
    .y     (_col_3_d_x4_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1308:100
    .z     (_col_3_n_u4_1_z)
  );
  ADD col_3_n_v4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1317:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_d_x8_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1315:100
    .y     (_delay_INT16_193_2304_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2322:118
    .z     (_col_3_n_v4_1_z)
  );
  SHR_3 col_3_n_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1318:83
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_v4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1317:100
    .z     (_col_3_n_x4_1_z)
  );
  dup_2 col_3_d_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1319:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1318:83
    .y     (_col_3_d_x4_1_y),
    .z     (_col_3_d_x4_1_z)
  );
  MUL col_3_n_u5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1320:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_w1_add_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1294:85
    .y     (_col_3_d_x5_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1309:100
    .z     (_col_3_n_u5_1_z)
  );
  SUB col_3_n_v5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1321:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_d_x8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1315:100
    .y     (_delay_INT16_178_1936_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1954:118
    .z     (_col_3_n_v5_1_z)
  );
  SHR_3 col_3_n_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1322:83
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_v5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1321:100
    .z     (_col_3_n_x5_1_z)
  );
  dup_2 col_3_d_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1323:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1322:83
    .y     (_col_3_d_x5_1_y),
    .z     (_col_3_d_x5_1_z)
  );
  ADD col_3_n_u8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1324:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_56_1935_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1953:114
    .y     (_col_3_d_x7_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1311:100
    .z     (_col_3_n_u8_1_z)
  );
  MUL col_3_n_v8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1325:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_w3_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1295:64
    .y     (_col_3_n_u8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1324:100
    .z     (_col_3_n_v8_1_z)
  );
  ADD col_3_n_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1326:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_v8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1325:100
    .y     (_col_3_n_c4_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1285:70
    .z     (_col_3_n_x8_1_z)
  );
  dup_2 col_3_d_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1327:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1326:100
    .y     (_col_3_d_x8_1_y),
    .z     (_col_3_d_x8_1_z)
  );
  MUL col_3_n_u6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1328:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_w3_sub_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1296:85
    .y     (_col_3_d_x6_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1310:100
    .z     (_col_3_n_u6_1_z)
  );
  SUB col_3_n_v6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1329:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_d_x8_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1327:100
    .y     (_delay_INT16_211_1934_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1952:118
    .z     (_col_3_n_v6_1_z)
  );
  SHR_3 col_3_n_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1330:83
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_v6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1329:100
    .z     (_col_3_n_x6_1_z)
  );
  dup_2 col_3_d_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1331:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1330:83
    .y     (_col_3_d_x6_1_y),
    .z     (_col_3_d_x6_1_z)
  );
  MUL col_3_n_u7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1332:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_w3_add_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1297:85
    .y     (_col_3_d_x7_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1311:100
    .z     (_col_3_n_u7_1_z)
  );
  SUB col_3_n_v7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1333:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_d_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1327:100
    .y     (_delay_INT16_176_1933_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1951:118
    .z     (_col_3_n_v7_1_z)
  );
  SHR_3 col_3_n_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1334:83
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_v7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1333:100
    .z     (_col_3_n_x7_1_z)
  );
  dup_2 col_3_d_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1335:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1334:83
    .y     (_col_3_d_x7_1_y),
    .z     (_col_3_d_x7_1_z)
  );
  ADD col_3_n_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1336:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_d_x0_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1304:100
    .y     (_delay_INT16_114_1932_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1950:118
    .z     (_col_3_n_x8_2_z)
  );
  dup_2 col_3_d_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1337:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1336:100
    .y     (_col_3_d_x8_2_y),
    .z     (_col_3_d_x8_2_z)
  );
  SUB col_3_n_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1338:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_d_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1304:100
    .y     (_delay_INT16_114_1931_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1949:118
    .z     (_col_3_n_x0_1_z)
  );
  dup_2 col_3_d_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1339:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1338:100
    .y     (_col_3_d_x0_1_y),
    .z     (_col_3_d_x0_1_z)
  );
  ADD col_3_n_u1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1340:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_d_x3_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1307:100
    .y     (_delay_INT16_133_2042_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2060:118
    .z     (_col_3_n_u1_1_z)
  );
  MUL col_3_n_v1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1341:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1298:64
    .y     (_col_3_n_u1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1340:100
    .z     (_col_3_n_v1_1_z)
  );
  ADD col_3_n_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1342:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_v1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1341:100
    .y     (_col_3_n_c4_2_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1286:70
    .z     (_col_3_n_x1_1_z)
  );
  dup_2 col_3_d_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1343:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1342:100
    .y     (_col_3_d_x1_1_y),
    .z     (_col_3_d_x1_1_z)
  );
  MUL col_3_n_u2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1344:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_w2_add_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1300:85
    .y     (_col_3_d_x2_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1306:100
    .z     (_col_3_n_u2_1_z)
  );
  SUB col_3_n_v2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1345:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_d_x1_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1343:100
    .y     (_delay_INT16_338_2013_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2031:118
    .z     (_col_3_n_v2_1_z)
  );
  SHR_3 col_3_n_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1346:83
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_v2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1345:100
    .z     (_col_3_n_x2_1_z)
  );
  dup_2 col_3_d_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1347:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1346:83
    .y     (_col_3_d_x2_1_y),
    .z     (_col_3_d_x2_1_z)
  );
  MUL col_3_n_u3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1348:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_w2_sub_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1299:85
    .y     (_col_3_d_x3_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1307:100
    .z     (_col_3_n_u3_1_z)
  );
  ADD col_3_n_v3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1349:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_d_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1343:100
    .y     (_delay_INT16_226_2322_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2340:118
    .z     (_col_3_n_v3_1_z)
  );
  SHR_3 col_3_n_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1350:83
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_v3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1349:100
    .z     (_col_3_n_x3_1_z)
  );
  dup_2 col_3_d_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1351:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1350:83
    .y     (_col_3_d_x3_1_y),
    .z     (_col_3_d_x3_1_z)
  );
  ADD col_3_n_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1352:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_d_x4_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1319:100
    .y     (_delay_INT16_1_1930_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1948:110
    .z     (_col_3_n_x1_2_z)
  );
  dup_2 col_3_d_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1353:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1352:100
    .y     (_col_3_d_x1_2_y),
    .z     (_col_3_d_x1_2_z)
  );
  SUB col_3_n_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1354:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_d_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1319:100
    .y     (_delay_INT16_1_1929_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1947:110
    .z     (_col_3_n_x4_2_z)
  );
  dup_2 col_3_d_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1355:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1354:100
    .y     (_col_3_d_x4_2_y),
    .z     (_col_3_d_x4_2_z)
  );
  ADD col_3_n_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1356:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_187_2051_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2069:118
    .y     (_col_3_d_x7_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1335:100
    .z     (_col_3_n_x6_2_z)
  );
  dup_2 col_3_d_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1357:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1356:100
    .y     (_col_3_d_x6_2_y),
    .z     (_col_3_d_x6_2_z)
  );
  SUB col_3_n_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1358:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_187_2225_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2243:118
    .y     (_col_3_d_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1335:100
    .z     (_col_3_n_x5_2_z)
  );
  dup_2 col_3_d_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1359:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1358:100
    .y     (_col_3_d_x5_2_y),
    .z     (_col_3_d_x5_2_z)
  );
  ADD col_3_n_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1360:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_59_1927_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1945:114
    .y     (_col_3_d_x3_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1351:100
    .z     (_col_3_n_x7_2_z)
  );
  dup_2 col_3_d_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1361:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1360:100
    .y     (_col_3_d_x7_2_y),
    .z     (_col_3_d_x7_2_z)
  );
  SUB col_3_n_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1362:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_59_1926_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1944:114
    .y     (_col_3_d_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1351:100
    .z     (_col_3_n_x8_3_z)
  );
  dup_2 col_3_d_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1363:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1362:100
    .y     (_col_3_d_x8_3_y),
    .z     (_col_3_d_x8_3_z)
  );
  ADD col_3_n_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1364:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_90_1925_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1943:114
    .y     (_col_3_d_x2_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1347:100
    .z     (_col_3_n_x3_2_z)
  );
  dup_2 col_3_d_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1365:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1364:100
    .y     (_col_3_d_x3_2_y),
    .z     (_col_3_d_x3_2_z)
  );
  SUB col_3_n_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1366:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_90_1924_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1942:114
    .y     (_col_3_d_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1347:100
    .z     (_col_3_n_x0_2_z)
  );
  dup_2 col_3_d_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1367:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1366:100
    .y     (_col_3_d_x0_2_y),
    .z     (_col_3_d_x0_2_z)
  );
  ADD col_3_n_u2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1368:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_140_1922_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1940:118
    .y     (_col_3_d_x5_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1359:100
    .z     (_col_3_n_u2_2_z)
  );
  MUL col_3_n_v2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1369:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_c181_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1289:76
    .y     (_col_3_n_u2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1368:100
    .z     (_col_3_n_v2_2_z)
  );
  ADD col_3_n_w2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1370:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_v2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1369:100
    .y     (_col_3_n_c128_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1287:76
    .z     (_col_3_n_w2_2_z)
  );
  SHR_8 col_3_n_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1371:83
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_w2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1370:100
    .z     (_col_3_n_x2_2_z)
  );
  dup_2 col_3_d_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1372:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1371:83
    .y     (_col_3_d_x2_2_y),
    .z     (_col_3_d_x2_2_z)
  );
  SUB col_3_n_u4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1373:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_140_1920_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1938:118
    .y     (_col_3_d_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1359:100
    .z     (_col_3_n_u4_3_z)
  );
  MUL col_3_n_v4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1374:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_c181_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1290:76
    .y     (_col_3_n_u4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1373:100
    .z     (_col_3_n_v4_3_z)
  );
  ADD col_3_n_w4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1375:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_v4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1374:100
    .y     (_col_3_n_c128_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1288:76
    .z     (_col_3_n_w4_3_z)
  );
  SHR_8 col_3_n_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1376:83
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_w4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1375:100
    .z     (_col_3_n_x4_3_z)
  );
  dup_2 col_3_d_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1377:100
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1376:83
    .y     (_col_3_d_x4_3_y),
    .z     (_col_3_d_x4_3_z)
  );
  ADD col_3_n_tmp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1378:105
    .clock (clock),
    .reset (reset),
    .x     (_col_3_d_x7_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1361:100
    .y     (_delay_INT16_99_1916_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1934:114
    .z     (_col_3_n_tmp_0_z)
  );
  SHR_14 col_3_n_val_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1379:87
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_tmp_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1378:105
    .z     (_col_3_n_val_0_z)
  );
  CLIP col_3_n_clp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1380:87
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_val_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1379:87
    .z     (n_out_0_3_x)
  );
  ADD col_3_n_tmp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1381:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_351_1915_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1933:118
    .y     (_col_3_d_x2_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1372:100
    .z     (_col_3_n_tmp_1_z)
  );
  SHR_14 col_3_n_val_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1382:87
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_tmp_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1381:105
    .z     (_col_3_n_val_1_z)
  );
  CLIP col_3_n_clp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1383:87
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_val_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1382:87
    .z     (n_out_1_3_x)
  );
  ADD col_3_n_tmp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1384:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_222_2115_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2133:118
    .y     (_col_3_d_x4_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1377:100
    .z     (_col_3_n_tmp_2_z)
  );
  SHR_14 col_3_n_val_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1385:87
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_tmp_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1384:105
    .z     (_col_3_n_val_2_z)
  );
  CLIP col_3_n_clp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1386:87
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_val_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1385:87
    .z     (n_out_2_3_x)
  );
  ADD col_3_n_tmp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1387:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_1_1914_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1932:110
    .y     (_col_3_d_x6_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1357:100
    .z     (_col_3_n_tmp_3_z)
  );
  SHR_14 col_3_n_val_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1388:87
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_tmp_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1387:105
    .z     (_col_3_n_val_3_z)
  );
  CLIP col_3_n_clp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1389:87
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_val_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1388:87
    .z     (n_out_3_3_x)
  );
  SUB col_3_n_tmp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1390:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_1_1913_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1931:110
    .y     (_col_3_d_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1357:100
    .z     (_col_3_n_tmp_4_z)
  );
  SHR_14 col_3_n_val_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1391:87
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_tmp_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1390:105
    .z     (_col_3_n_val_4_z)
  );
  CLIP col_3_n_clp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1392:87
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_val_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1391:87
    .z     (n_out_4_3_x)
  );
  SUB col_3_n_tmp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1393:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_222_1912_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1930:118
    .y     (_col_3_d_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1377:100
    .z     (_col_3_n_tmp_5_z)
  );
  SHR_14 col_3_n_val_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1394:87
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_tmp_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1393:105
    .z     (_col_3_n_val_5_z)
  );
  CLIP col_3_n_clp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1395:87
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_val_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1394:87
    .z     (n_out_5_3_x)
  );
  SUB col_3_n_tmp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1396:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_351_1911_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1929:118
    .y     (_col_3_d_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1372:100
    .z     (_col_3_n_tmp_6_z)
  );
  SHR_14 col_3_n_val_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1397:87
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_tmp_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1396:105
    .z     (_col_3_n_val_6_z)
  );
  CLIP col_3_n_clp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1398:87
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_val_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1397:87
    .z     (n_out_6_3_x)
  );
  SUB col_3_n_tmp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1399:105
    .clock (clock),
    .reset (reset),
    .x     (_col_3_d_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1361:100
    .y     (_delay_INT16_99_2073_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2091:114
    .z     (_col_3_n_tmp_7_z)
  );
  SHR_14 col_3_n_val_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1400:87
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_tmp_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1399:105
    .z     (_col_3_n_val_7_z)
  );
  CLIP col_3_n_clp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1401:87
    .clock (clock),
    .reset (reset),
    .x     (_col_3_n_val_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1400:87
    .z     (n_out_7_3_x)
  );
  C4 col_4_n_c4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1402:70
    .clock (clock),
    .reset (reset),
    .value (_col_4_n_c4_0_value)
  );
  C4 col_4_n_c4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1403:70
    .clock (clock),
    .reset (reset),
    .value (_col_4_n_c4_1_value)
  );
  C4 col_4_n_c4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1404:70
    .clock (clock),
    .reset (reset),
    .value (_col_4_n_c4_2_value)
  );
  C128 col_4_n_c128_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1405:76
    .clock (clock),
    .reset (reset),
    .value (_col_4_n_c128_0_value)
  );
  C128 col_4_n_c128_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1406:76
    .clock (clock),
    .reset (reset),
    .value (_col_4_n_c128_1_value)
  );
  C181 col_4_n_c181_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1407:76
    .clock (clock),
    .reset (reset),
    .value (_col_4_n_c181_0_value)
  );
  C181 col_4_n_c181_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1408:76
    .clock (clock),
    .reset (reset),
    .value (_col_4_n_c181_1_value)
  );
  C8192 col_4_n_c8192 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1409:73
    .clock (clock),
    .reset (reset),
    .value (_col_4_n_c8192_value)
  );
  W7 col_4_n_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1410:64
    .clock (clock),
    .reset (reset),
    .value (_col_4_n_w7_value)
  );
  W1_sub_W7 col_4_n_w1_sub_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1411:85
    .clock (clock),
    .reset (reset),
    .value (_col_4_n_w1_sub_w7_value)
  );
  W1_add_W7 col_4_n_w1_add_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1412:85
    .clock (clock),
    .reset (reset),
    .value (_col_4_n_w1_add_w7_value)
  );
  W3 col_4_n_w3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1413:64
    .clock (clock),
    .reset (reset),
    .value (_col_4_n_w3_value)
  );
  W3_sub_W5 col_4_n_w3_sub_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1414:85
    .clock (clock),
    .reset (reset),
    .value (_col_4_n_w3_sub_w5_value)
  );
  W3_add_W5 col_4_n_w3_add_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1415:85
    .clock (clock),
    .reset (reset),
    .value (_col_4_n_w3_add_w5_value)
  );
  W6 col_4_n_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1416:64
    .clock (clock),
    .reset (reset),
    .value (_col_4_n_w6_value)
  );
  W2_sub_W6 col_4_n_w2_sub_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1417:85
    .clock (clock),
    .reset (reset),
    .value (_col_4_n_w2_sub_w6_value)
  );
  W2_add_W6 col_4_n_w2_add_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1418:85
    .clock (clock),
    .reset (reset),
    .value (_col_4_n_w2_add_w6_value)
  );
  SHL_8 col_4_n_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1419:83
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_shr_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:629:87
    .z     (_col_4_n_x1_0_z)
  );
  SHL_8 col_4_n_t0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1420:83
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_shr_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:237:87
    .z     (_col_4_n_t0_0_z)
  );
  ADD col_4_n_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1421:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_t0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1420:83
    .y     (_col_4_n_c8192_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1409:73
    .z     (_col_4_n_x0_0_z)
  );
  dup_2 col_4_d_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1422:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1421:100
    .y     (_col_4_d_x0_0_y),
    .z     (_col_4_d_x0_0_z)
  );
  dup_2 col_4_d_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1423:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1419:83
    .y     (_col_4_d_x1_0_y),
    .z     (_col_4_d_x1_0_z)
  );
  dup_2 col_4_d_x2_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1424:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_shr_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:825:87
    .y     (_col_4_d_x2_0_y),
    .z     (_col_4_d_x2_0_z)
  );
  dup_2 col_4_d_x3_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1425:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_shr_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:433:87
    .y     (_col_4_d_x3_0_y),
    .z     (_col_4_d_x3_0_z)
  );
  dup_2 col_4_d_x4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1426:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_shr_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:335:87
    .y     (_col_4_d_x4_0_y),
    .z     (_col_4_d_x4_0_z)
  );
  dup_2 col_4_d_x5_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1427:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_shr_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:923:87
    .y     (_col_4_d_x5_0_y),
    .z     (_col_4_d_x5_0_z)
  );
  dup_2 col_4_d_x6_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1428:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_shr_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:727:87
    .y     (_col_4_d_x6_0_y),
    .z     (_col_4_d_x6_0_z)
  );
  dup_2 col_4_d_x7_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1429:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_shr_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:531:87
    .y     (_col_4_d_x7_0_y),
    .z     (_col_4_d_x7_0_z)
  );
  ADD col_4_n_u8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1430:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x4_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1426:100
    .y     (_delay_INT16_6_2321_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2339:110
    .z     (_col_4_n_u8_0_z)
  );
  MUL col_4_n_v8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1431:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1410:64
    .y     (_col_4_n_u8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1430:100
    .z     (_col_4_n_v8_0_z)
  );
  ADD col_4_n_x8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1432:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_v8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1431:100
    .y     (_col_4_n_c4_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1402:70
    .z     (_col_4_n_x8_0_z)
  );
  dup_2 col_4_d_x8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1433:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1432:100
    .y     (_col_4_d_x8_0_y),
    .z     (_col_4_d_x8_0_z)
  );
  MUL col_4_n_u4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1434:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_w1_sub_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1411:85
    .y     (_col_4_d_x4_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1426:100
    .z     (_col_4_n_u4_1_z)
  );
  ADD col_4_n_v4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1435:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x8_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1433:100
    .y     (_delay_INT16_231_1928_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1946:118
    .z     (_col_4_n_v4_1_z)
  );
  SHR_3 col_4_n_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1436:83
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_v4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1435:100
    .z     (_col_4_n_x4_1_z)
  );
  dup_2 col_4_d_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1437:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1436:83
    .y     (_col_4_d_x4_1_y),
    .z     (_col_4_d_x4_1_z)
  );
  MUL col_4_n_u5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1438:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_w1_add_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1412:85
    .y     (_col_4_d_x5_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1427:100
    .z     (_col_4_n_u5_1_z)
  );
  SUB col_4_n_v5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1439:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1433:100
    .y     (_delay_INT16_235_2224_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2242:118
    .z     (_col_4_n_v5_1_z)
  );
  SHR_3 col_4_n_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1440:83
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_v5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1439:100
    .z     (_col_4_n_x5_1_z)
  );
  dup_2 col_4_d_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1441:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1440:83
    .y     (_col_4_d_x5_1_y),
    .z     (_col_4_d_x5_1_z)
  );
  ADD col_4_n_u8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1442:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x6_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1428:100
    .y     (_delay_INT16_100_2230_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2248:118
    .z     (_col_4_n_u8_1_z)
  );
  MUL col_4_n_v8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1443:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_w3_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1413:64
    .y     (_col_4_n_u8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1442:100
    .z     (_col_4_n_v8_1_z)
  );
  ADD col_4_n_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1444:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_v8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1443:100
    .y     (_col_4_n_c4_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1403:70
    .z     (_col_4_n_x8_1_z)
  );
  dup_2 col_4_d_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1445:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1444:100
    .y     (_col_4_d_x8_1_y),
    .z     (_col_4_d_x8_1_z)
  );
  MUL col_4_n_u6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1446:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_w3_sub_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1414:85
    .y     (_col_4_d_x6_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1428:100
    .z     (_col_4_n_u6_1_z)
  );
  SUB col_4_n_v6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1447:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x8_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1445:100
    .y     (_delay_INT16_7_1923_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1941:110
    .z     (_col_4_n_v6_1_z)
  );
  SHR_3 col_4_n_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1448:83
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_v6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1447:100
    .z     (_col_4_n_x6_1_z)
  );
  dup_2 col_4_d_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1449:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1448:83
    .y     (_col_4_d_x6_1_y),
    .z     (_col_4_d_x6_1_z)
  );
  MUL col_4_n_u7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1450:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_w3_add_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1415:85
    .y     (_col_4_d_x7_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1429:100
    .z     (_col_4_n_u7_1_z)
  );
  SUB col_4_n_v7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1451:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1445:100
    .y     (_delay_INT16_106_1921_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1939:118
    .z     (_col_4_n_v7_1_z)
  );
  SHR_3 col_4_n_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1452:83
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_v7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1451:100
    .z     (_col_4_n_x7_1_z)
  );
  dup_2 col_4_d_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1453:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1452:83
    .y     (_col_4_d_x7_1_y),
    .z     (_col_4_d_x7_1_z)
  );
  ADD col_4_n_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1454:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_125_1919_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1937:118
    .y     (_col_4_d_x1_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1423:100
    .z     (_col_4_n_x8_2_z)
  );
  dup_2 col_4_d_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1455:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1454:100
    .y     (_col_4_d_x8_2_y),
    .z     (_col_4_d_x8_2_z)
  );
  SUB col_4_n_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1456:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_125_1918_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1936:118
    .y     (_col_4_d_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1423:100
    .z     (_col_4_n_x0_1_z)
  );
  dup_2 col_4_d_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1457:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1456:100
    .y     (_col_4_d_x0_1_y),
    .z     (_col_4_d_x0_1_z)
  );
  ADD col_4_n_u1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1458:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x3_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1425:100
    .y     (_delay_INT16_27_1917_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1935:114
    .z     (_col_4_n_u1_1_z)
  );
  MUL col_4_n_v1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1459:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1416:64
    .y     (_col_4_n_u1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1458:100
    .z     (_col_4_n_v1_1_z)
  );
  ADD col_4_n_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1460:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_v1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1459:100
    .y     (_col_4_n_c4_2_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1404:70
    .z     (_col_4_n_x1_1_z)
  );
  dup_2 col_4_d_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1461:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1460:100
    .y     (_col_4_d_x1_1_y),
    .z     (_col_4_d_x1_1_z)
  );
  MUL col_4_n_u2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1462:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_w2_add_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1418:85
    .y     (_col_4_d_x2_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1424:100
    .z     (_col_4_n_u2_1_z)
  );
  SUB col_4_n_v2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1463:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x1_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1461:100
    .y     (_delay_INT16_207_1910_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1928:118
    .z     (_col_4_n_v2_1_z)
  );
  SHR_3 col_4_n_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1464:83
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_v2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1463:100
    .z     (_col_4_n_x2_1_z)
  );
  dup_2 col_4_d_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1465:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1464:83
    .y     (_col_4_d_x2_1_y),
    .z     (_col_4_d_x2_1_z)
  );
  MUL col_4_n_u3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1466:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_w2_sub_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1417:85
    .y     (_col_4_d_x3_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1425:100
    .z     (_col_4_n_u3_1_z)
  );
  ADD col_4_n_v3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1467:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1461:100
    .y     (_delay_INT16_159_1909_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1927:118
    .z     (_col_4_n_v3_1_z)
  );
  SHR_3 col_4_n_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1468:83
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_v3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1467:100
    .z     (_col_4_n_x3_1_z)
  );
  dup_2 col_4_d_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1469:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1468:83
    .y     (_col_4_d_x3_1_y),
    .z     (_col_4_d_x3_1_z)
  );
  ADD col_4_n_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1470:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x4_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1437:100
    .y     (_delay_INT16_131_2083_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2101:118
    .z     (_col_4_n_x1_2_z)
  );
  dup_2 col_4_d_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1471:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1470:100
    .y     (_col_4_d_x1_2_y),
    .z     (_col_4_d_x1_2_z)
  );
  SUB col_4_n_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1472:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1437:100
    .y     (_delay_INT16_131_1908_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1926:118
    .z     (_col_4_n_x4_2_z)
  );
  dup_2 col_4_d_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1473:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1472:100
    .y     (_col_4_d_x4_2_y),
    .z     (_col_4_d_x4_2_z)
  );
  ADD col_4_n_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1474:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x5_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1441:100
    .y     (_delay_INT16_165_1907_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1925:118
    .z     (_col_4_n_x6_2_z)
  );
  dup_2 col_4_d_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1475:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1474:100
    .y     (_col_4_d_x6_2_y),
    .z     (_col_4_d_x6_2_z)
  );
  SUB col_4_n_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1476:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1441:100
    .y     (_delay_INT16_165_1906_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1924:118
    .z     (_col_4_n_x5_2_z)
  );
  dup_2 col_4_d_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1477:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1476:100
    .y     (_col_4_d_x5_2_y),
    .z     (_col_4_d_x5_2_z)
  );
  ADD col_4_n_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1478:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_21_1905_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1923:114
    .y     (_col_4_d_x3_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1469:100
    .z     (_col_4_n_x7_2_z)
  );
  dup_2 col_4_d_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1479:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1478:100
    .y     (_col_4_d_x7_2_y),
    .z     (_col_4_d_x7_2_z)
  );
  SUB col_4_n_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1480:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_21_2005_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2023:114
    .y     (_col_4_d_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1469:100
    .z     (_col_4_n_x8_3_z)
  );
  dup_2 col_4_d_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1481:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1480:100
    .y     (_col_4_d_x8_3_y),
    .z     (_col_4_d_x8_3_z)
  );
  ADD col_4_n_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1482:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x0_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1457:100
    .y     (_delay_INT16_17_1967_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1985:114
    .z     (_col_4_n_x3_2_z)
  );
  dup_2 col_4_d_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1483:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1482:100
    .y     (_col_4_d_x3_2_y),
    .z     (_col_4_d_x3_2_z)
  );
  SUB col_4_n_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1484:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1457:100
    .y     (_delay_INT16_17_1904_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1922:114
    .z     (_col_4_n_x0_2_z)
  );
  dup_2 col_4_d_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1485:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1484:100
    .y     (_col_4_d_x0_2_y),
    .z     (_col_4_d_x0_2_z)
  );
  ADD col_4_n_u2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1486:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x4_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1473:100
    .y     (_col_4_d_x5_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1477:100
    .z     (_col_4_n_u2_2_z)
  );
  MUL col_4_n_v2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1487:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_c181_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1407:76
    .y     (_col_4_n_u2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1486:100
    .z     (_col_4_n_v2_2_z)
  );
  ADD col_4_n_w2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1488:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_v2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1487:100
    .y     (_col_4_n_c128_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1405:76
    .z     (_col_4_n_w2_2_z)
  );
  SHR_8 col_4_n_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1489:83
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_w2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1488:100
    .z     (_col_4_n_x2_2_z)
  );
  dup_2 col_4_d_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1490:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1489:83
    .y     (_col_4_d_x2_2_y),
    .z     (_col_4_d_x2_2_z)
  );
  SUB col_4_n_u4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1491:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1473:100
    .y     (_col_4_d_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1477:100
    .z     (_col_4_n_u4_3_z)
  );
  MUL col_4_n_v4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1492:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_c181_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1408:76
    .y     (_col_4_n_u4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1491:100
    .z     (_col_4_n_v4_3_z)
  );
  ADD col_4_n_w4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1493:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_v4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1492:100
    .y     (_col_4_n_c128_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1406:76
    .z     (_col_4_n_w4_3_z)
  );
  SHR_8 col_4_n_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1494:83
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_w4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1493:100
    .z     (_col_4_n_x4_3_z)
  );
  dup_2 col_4_d_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1495:100
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1494:83
    .y     (_col_4_d_x4_3_y),
    .z     (_col_4_d_x4_3_z)
  );
  ADD col_4_n_tmp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1496:105
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x7_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1479:100
    .y     (_delay_INT16_38_1903_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1921:114
    .z     (_col_4_n_tmp_0_z)
  );
  SHR_14 col_4_n_val_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1497:87
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_tmp_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1496:105
    .z     (_col_4_n_val_0_z)
  );
  CLIP col_4_n_clp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1498:87
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_val_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1497:87
    .z     (n_out_0_4_x)
  );
  ADD col_4_n_tmp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1499:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_119_2313_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2331:118
    .y     (_col_4_d_x2_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1490:100
    .z     (_col_4_n_tmp_1_z)
  );
  SHR_14 col_4_n_val_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1500:87
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_tmp_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1499:105
    .z     (_col_4_n_val_1_z)
  );
  CLIP col_4_n_clp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1501:87
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_val_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1500:87
    .z     (n_out_1_4_x)
  );
  ADD col_4_n_tmp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1502:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_334_1902_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1920:118
    .y     (_col_4_d_x4_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1495:100
    .z     (_col_4_n_tmp_2_z)
  );
  SHR_14 col_4_n_val_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1503:87
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_tmp_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1502:105
    .z     (_col_4_n_val_2_z)
  );
  CLIP col_4_n_clp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1504:87
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_val_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1503:87
    .z     (n_out_2_4_x)
  );
  ADD col_4_n_tmp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1505:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_2_2058_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2076:110
    .y     (_col_4_d_x6_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1475:100
    .z     (_col_4_n_tmp_3_z)
  );
  SHR_14 col_4_n_val_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1506:87
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_tmp_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1505:105
    .z     (_col_4_n_val_3_z)
  );
  CLIP col_4_n_clp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1507:87
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_val_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1506:87
    .z     (n_out_3_4_x)
  );
  SUB col_4_n_tmp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1508:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_2_1901_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1919:110
    .y     (_col_4_d_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1475:100
    .z     (_col_4_n_tmp_4_z)
  );
  SHR_14 col_4_n_val_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1509:87
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_tmp_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1508:105
    .z     (_col_4_n_val_4_z)
  );
  CLIP col_4_n_clp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1510:87
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_val_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1509:87
    .z     (n_out_4_4_x)
  );
  SUB col_4_n_tmp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1511:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_334_1900_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1918:118
    .y     (_col_4_d_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1495:100
    .z     (_col_4_n_tmp_5_z)
  );
  SHR_14 col_4_n_val_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1512:87
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_tmp_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1511:105
    .z     (_col_4_n_val_5_z)
  );
  CLIP col_4_n_clp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1513:87
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_val_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1512:87
    .z     (n_out_5_4_x)
  );
  SUB col_4_n_tmp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1514:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_119_2158_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2176:118
    .y     (_col_4_d_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1490:100
    .z     (_col_4_n_tmp_6_z)
  );
  SHR_14 col_4_n_val_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1515:87
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_tmp_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1514:105
    .z     (_col_4_n_val_6_z)
  );
  CLIP col_4_n_clp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1516:87
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_val_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1515:87
    .z     (n_out_6_4_x)
  );
  SUB col_4_n_tmp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1517:105
    .clock (clock),
    .reset (reset),
    .x     (_col_4_d_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1479:100
    .y     (_delay_INT16_38_2025_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2043:114
    .z     (_col_4_n_tmp_7_z)
  );
  SHR_14 col_4_n_val_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1518:87
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_tmp_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1517:105
    .z     (_col_4_n_val_7_z)
  );
  CLIP col_4_n_clp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1519:87
    .clock (clock),
    .reset (reset),
    .x     (_col_4_n_val_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1518:87
    .z     (n_out_7_4_x)
  );
  C4 col_5_n_c4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1520:70
    .clock (clock),
    .reset (reset),
    .value (_col_5_n_c4_0_value)
  );
  C4 col_5_n_c4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1521:70
    .clock (clock),
    .reset (reset),
    .value (_col_5_n_c4_1_value)
  );
  C4 col_5_n_c4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1522:70
    .clock (clock),
    .reset (reset),
    .value (_col_5_n_c4_2_value)
  );
  C128 col_5_n_c128_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1523:76
    .clock (clock),
    .reset (reset),
    .value (_col_5_n_c128_0_value)
  );
  C128 col_5_n_c128_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1524:76
    .clock (clock),
    .reset (reset),
    .value (_col_5_n_c128_1_value)
  );
  C181 col_5_n_c181_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1525:76
    .clock (clock),
    .reset (reset),
    .value (_col_5_n_c181_0_value)
  );
  C181 col_5_n_c181_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1526:76
    .clock (clock),
    .reset (reset),
    .value (_col_5_n_c181_1_value)
  );
  C8192 col_5_n_c8192 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1527:73
    .clock (clock),
    .reset (reset),
    .value (_col_5_n_c8192_value)
  );
  W7 col_5_n_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1528:64
    .clock (clock),
    .reset (reset),
    .value (_col_5_n_w7_value)
  );
  W1_sub_W7 col_5_n_w1_sub_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1529:85
    .clock (clock),
    .reset (reset),
    .value (_col_5_n_w1_sub_w7_value)
  );
  W1_add_W7 col_5_n_w1_add_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1530:85
    .clock (clock),
    .reset (reset),
    .value (_col_5_n_w1_add_w7_value)
  );
  W3 col_5_n_w3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1531:64
    .clock (clock),
    .reset (reset),
    .value (_col_5_n_w3_value)
  );
  W3_sub_W5 col_5_n_w3_sub_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1532:85
    .clock (clock),
    .reset (reset),
    .value (_col_5_n_w3_sub_w5_value)
  );
  W3_add_W5 col_5_n_w3_add_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1533:85
    .clock (clock),
    .reset (reset),
    .value (_col_5_n_w3_add_w5_value)
  );
  W6 col_5_n_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1534:64
    .clock (clock),
    .reset (reset),
    .value (_col_5_n_w6_value)
  );
  W2_sub_W6 col_5_n_w2_sub_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1535:85
    .clock (clock),
    .reset (reset),
    .value (_col_5_n_w2_sub_w6_value)
  );
  W2_add_W6 col_5_n_w2_add_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1536:85
    .clock (clock),
    .reset (reset),
    .value (_col_5_n_w2_add_w6_value)
  );
  SHL_8 col_5_n_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1537:83
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_shr_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:631:87
    .z     (_col_5_n_x1_0_z)
  );
  SHL_8 col_5_n_t0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1538:83
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_shr_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:239:87
    .z     (_col_5_n_t0_0_z)
  );
  ADD col_5_n_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1539:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_t0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1538:83
    .y     (_col_5_n_c8192_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1527:73
    .z     (_col_5_n_x0_0_z)
  );
  dup_2 col_5_d_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1540:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1539:100
    .y     (_col_5_d_x0_0_y),
    .z     (_col_5_d_x0_0_z)
  );
  dup_2 col_5_d_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1541:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1537:83
    .y     (_col_5_d_x1_0_y),
    .z     (_col_5_d_x1_0_z)
  );
  dup_2 col_5_d_x2_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1542:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_shr_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:827:87
    .y     (_col_5_d_x2_0_y),
    .z     (_col_5_d_x2_0_z)
  );
  dup_2 col_5_d_x3_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1543:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_shr_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:435:87
    .y     (_col_5_d_x3_0_y),
    .z     (_col_5_d_x3_0_z)
  );
  dup_2 col_5_d_x4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1544:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_shr_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:337:87
    .y     (_col_5_d_x4_0_y),
    .z     (_col_5_d_x4_0_z)
  );
  dup_2 col_5_d_x5_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1545:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_shr_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:925:87
    .y     (_col_5_d_x5_0_y),
    .z     (_col_5_d_x5_0_z)
  );
  dup_2 col_5_d_x6_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1546:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_shr_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:729:87
    .y     (_col_5_d_x6_0_y),
    .z     (_col_5_d_x6_0_z)
  );
  dup_2 col_5_d_x7_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1547:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_shr_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:533:87
    .y     (_col_5_d_x7_0_y),
    .z     (_col_5_d_x7_0_z)
  );
  ADD col_5_n_u8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1548:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_d_x4_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1544:100
    .y     (_delay_INT16_26_1899_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1917:114
    .z     (_col_5_n_u8_0_z)
  );
  MUL col_5_n_v8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1549:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1528:64
    .y     (_col_5_n_u8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1548:100
    .z     (_col_5_n_v8_0_z)
  );
  ADD col_5_n_x8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1550:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_v8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1549:100
    .y     (_col_5_n_c4_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1520:70
    .z     (_col_5_n_x8_0_z)
  );
  dup_2 col_5_d_x8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1551:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1550:100
    .y     (_col_5_d_x8_0_y),
    .z     (_col_5_d_x8_0_z)
  );
  MUL col_5_n_u4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1552:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_w1_sub_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1529:85
    .y     (_col_5_d_x4_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1544:100
    .z     (_col_5_n_u4_1_z)
  );
  ADD col_5_n_v4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1553:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_6_1898_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1916:110
    .y     (_col_5_n_u4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1552:100
    .z     (_col_5_n_v4_1_z)
  );
  SHR_3 col_5_n_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1554:83
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_v4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1553:100
    .z     (_col_5_n_x4_1_z)
  );
  dup_2 col_5_d_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1555:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1554:83
    .y     (_col_5_d_x4_1_y),
    .z     (_col_5_d_x4_1_z)
  );
  MUL col_5_n_u5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1556:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_w1_add_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1530:85
    .y     (_col_5_d_x5_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1545:100
    .z     (_col_5_n_u5_1_z)
  );
  SUB col_5_n_v5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1557:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_d_x8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1551:100
    .y     (_delay_INT16_14_1897_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1915:114
    .z     (_col_5_n_v5_1_z)
  );
  SHR_3 col_5_n_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1558:83
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_v5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1557:100
    .z     (_col_5_n_x5_1_z)
  );
  dup_2 col_5_d_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1559:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1558:83
    .y     (_col_5_d_x5_1_y),
    .z     (_col_5_d_x5_1_z)
  );
  ADD col_5_n_u8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1560:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_82_2138_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2156:114
    .y     (_col_5_d_x7_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1547:100
    .z     (_col_5_n_u8_1_z)
  );
  MUL col_5_n_v8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1561:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_w3_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1531:64
    .y     (_col_5_n_u8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1560:100
    .z     (_col_5_n_v8_1_z)
  );
  ADD col_5_n_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1562:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_v8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1561:100
    .y     (_col_5_n_c4_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1521:70
    .z     (_col_5_n_x8_1_z)
  );
  dup_2 col_5_d_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1563:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1562:100
    .y     (_col_5_d_x8_1_y),
    .z     (_col_5_d_x8_1_z)
  );
  MUL col_5_n_u6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1564:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_w3_sub_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1532:85
    .y     (_col_5_d_x6_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1546:100
    .z     (_col_5_n_u6_1_z)
  );
  SUB col_5_n_v6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1565:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_d_x8_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1563:100
    .y     (_delay_INT16_230_1896_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1914:118
    .z     (_col_5_n_v6_1_z)
  );
  SHR_3 col_5_n_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1566:83
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_v6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1565:100
    .z     (_col_5_n_x6_1_z)
  );
  dup_2 col_5_d_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1567:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1566:83
    .y     (_col_5_d_x6_1_y),
    .z     (_col_5_d_x6_1_z)
  );
  MUL col_5_n_u7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1568:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_w3_add_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1533:85
    .y     (_col_5_d_x7_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1547:100
    .z     (_col_5_n_u7_1_z)
  );
  SUB col_5_n_v7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1569:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_d_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1563:100
    .y     (_delay_INT16_130_1895_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1913:118
    .z     (_col_5_n_v7_1_z)
  );
  SHR_3 col_5_n_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1570:83
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_v7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1569:100
    .z     (_col_5_n_x7_1_z)
  );
  dup_2 col_5_d_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1571:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1570:83
    .y     (_col_5_d_x7_1_y),
    .z     (_col_5_d_x7_1_z)
  );
  ADD col_5_n_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1572:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_121_1894_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1912:118
    .y     (_col_5_d_x1_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1541:100
    .z     (_col_5_n_x8_2_z)
  );
  dup_2 col_5_d_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1573:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1572:100
    .y     (_col_5_d_x8_2_y),
    .z     (_col_5_d_x8_2_z)
  );
  SUB col_5_n_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1574:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_121_2319_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2337:118
    .y     (_col_5_d_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1541:100
    .z     (_col_5_n_x0_1_z)
  );
  dup_2 col_5_d_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1575:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1574:100
    .y     (_col_5_d_x0_1_y),
    .z     (_col_5_d_x0_1_z)
  );
  ADD col_5_n_u1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1576:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_81_1893_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1911:114
    .y     (_col_5_d_x2_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1542:100
    .z     (_col_5_n_u1_1_z)
  );
  MUL col_5_n_v1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1577:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1534:64
    .y     (_col_5_n_u1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1576:100
    .z     (_col_5_n_v1_1_z)
  );
  ADD col_5_n_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1578:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_v1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1577:100
    .y     (_col_5_n_c4_2_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1522:70
    .z     (_col_5_n_x1_1_z)
  );
  dup_2 col_5_d_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1579:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1578:100
    .y     (_col_5_d_x1_1_y),
    .z     (_col_5_d_x1_1_z)
  );
  MUL col_5_n_u2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1580:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_w2_add_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1536:85
    .y     (_col_5_d_x2_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1542:100
    .z     (_col_5_n_u2_1_z)
  );
  SUB col_5_n_v2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1581:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_d_x1_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1579:100
    .y     (_delay_INT16_126_1892_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1910:118
    .z     (_col_5_n_v2_1_z)
  );
  SHR_3 col_5_n_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1582:83
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_v2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1581:100
    .z     (_col_5_n_x2_1_z)
  );
  dup_2 col_5_d_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1583:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1582:83
    .y     (_col_5_d_x2_1_y),
    .z     (_col_5_d_x2_1_z)
  );
  MUL col_5_n_u3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1584:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_w2_sub_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1535:85
    .y     (_col_5_d_x3_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1543:100
    .z     (_col_5_n_u3_1_z)
  );
  ADD col_5_n_v3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1585:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_d_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1579:100
    .y     (_delay_INT16_225_2177_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2195:118
    .z     (_col_5_n_v3_1_z)
  );
  SHR_3 col_5_n_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1586:83
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_v3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1585:100
    .z     (_col_5_n_x3_1_z)
  );
  dup_2 col_5_d_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1587:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1586:83
    .y     (_col_5_d_x3_1_y),
    .z     (_col_5_d_x3_1_z)
  );
  ADD col_5_n_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1588:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_378_2220_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2238:118
    .y     (_col_5_d_x6_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1567:100
    .z     (_col_5_n_x1_2_z)
  );
  dup_2 col_5_d_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1589:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1588:100
    .y     (_col_5_d_x1_2_y),
    .z     (_col_5_d_x1_2_z)
  );
  SUB col_5_n_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1590:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_378_1891_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1909:118
    .y     (_col_5_d_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1567:100
    .z     (_col_5_n_x4_2_z)
  );
  dup_2 col_5_d_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1591:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1590:100
    .y     (_col_5_d_x4_2_y),
    .z     (_col_5_d_x4_2_z)
  );
  ADD col_5_n_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1592:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_378_1947_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1965:118
    .y     (_col_5_d_x7_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1571:100
    .z     (_col_5_n_x6_2_z)
  );
  dup_2 col_5_d_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1593:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1592:100
    .y     (_col_5_d_x6_2_y),
    .z     (_col_5_d_x6_2_z)
  );
  SUB col_5_n_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1594:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_378_2314_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2332:118
    .y     (_col_5_d_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1571:100
    .z     (_col_5_n_x5_2_z)
  );
  dup_2 col_5_d_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1595:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1594:100
    .y     (_col_5_d_x5_2_y),
    .z     (_col_5_d_x5_2_z)
  );
  ADD col_5_n_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1596:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_61_2300_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2318:114
    .y     (_col_5_d_x3_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1587:100
    .z     (_col_5_n_x7_2_z)
  );
  dup_2 col_5_d_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1597:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1596:100
    .y     (_col_5_d_x7_2_y),
    .z     (_col_5_d_x7_2_z)
  );
  SUB col_5_n_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1598:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_61_2201_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2219:114
    .y     (_col_5_d_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1587:100
    .z     (_col_5_n_x8_3_z)
  );
  dup_2 col_5_d_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1599:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1598:100
    .y     (_col_5_d_x8_3_y),
    .z     (_col_5_d_x8_3_z)
  );
  ADD col_5_n_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1600:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_186_2193_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2211:118
    .y     (_col_5_d_x2_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1583:100
    .z     (_col_5_n_x3_2_z)
  );
  dup_2 col_5_d_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1601:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1600:100
    .y     (_col_5_d_x3_2_y),
    .z     (_col_5_d_x3_2_z)
  );
  SUB col_5_n_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1602:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_186_1890_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1908:118
    .y     (_col_5_d_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1583:100
    .z     (_col_5_n_x0_2_z)
  );
  dup_2 col_5_d_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1603:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1602:100
    .y     (_col_5_d_x0_2_y),
    .z     (_col_5_d_x0_2_z)
  );
  ADD col_5_n_u2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1604:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_d_x4_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1591:100
    .y     (_delay_INT16_24_2082_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2100:114
    .z     (_col_5_n_u2_2_z)
  );
  MUL col_5_n_v2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1605:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_c181_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1525:76
    .y     (_col_5_n_u2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1604:100
    .z     (_col_5_n_v2_2_z)
  );
  ADD col_5_n_w2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1606:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_v2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1605:100
    .y     (_col_5_n_c128_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1523:76
    .z     (_col_5_n_w2_2_z)
  );
  SHR_8 col_5_n_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1607:83
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_w2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1606:100
    .z     (_col_5_n_x2_2_z)
  );
  dup_2 col_5_d_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1608:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1607:83
    .y     (_col_5_d_x2_2_y),
    .z     (_col_5_d_x2_2_z)
  );
  SUB col_5_n_u4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1609:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_d_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1591:100
    .y     (_delay_INT16_24_2097_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2115:114
    .z     (_col_5_n_u4_3_z)
  );
  MUL col_5_n_v4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1610:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_c181_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1526:76
    .y     (_col_5_n_u4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1609:100
    .z     (_col_5_n_v4_3_z)
  );
  ADD col_5_n_w4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1611:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_v4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1610:100
    .y     (_col_5_n_c128_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1524:76
    .z     (_col_5_n_w4_3_z)
  );
  SHR_8 col_5_n_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1612:83
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_w4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1611:100
    .z     (_col_5_n_x4_3_z)
  );
  dup_2 col_5_d_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1613:100
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1612:83
    .y     (_col_5_d_x4_3_y),
    .z     (_col_5_d_x4_3_z)
  );
  ADD col_5_n_tmp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1614:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_80_2165_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2183:114
    .y     (_col_5_d_x1_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1589:100
    .z     (_col_5_n_tmp_0_z)
  );
  SHR_14 col_5_n_val_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1615:87
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_tmp_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1614:105
    .z     (_col_5_n_val_0_z)
  );
  CLIP col_5_n_clp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1616:87
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_val_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1615:87
    .z     (n_out_0_5_x)
  );
  ADD col_5_n_tmp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1617:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_180_2305_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2323:118
    .y     (_col_5_d_x2_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1608:100
    .z     (_col_5_n_tmp_1_z)
  );
  SHR_14 col_5_n_val_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1618:87
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_tmp_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1617:105
    .z     (_col_5_n_val_1_z)
  );
  CLIP col_5_n_clp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1619:87
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_val_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1618:87
    .z     (n_out_1_5_x)
  );
  ADD col_5_n_tmp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1620:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_288_2034_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2052:118
    .y     (_col_5_d_x4_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1613:100
    .z     (_col_5_n_tmp_2_z)
  );
  SHR_14 col_5_n_val_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1621:87
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_tmp_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1620:105
    .z     (_col_5_n_val_2_z)
  );
  CLIP col_5_n_clp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1622:87
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_val_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1621:87
    .z     (n_out_2_5_x)
  );
  ADD col_5_n_tmp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1623:105
    .clock (clock),
    .reset (reset),
    .x     (_col_5_d_x8_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1599:100
    .y     (_delay_INT16_57_1889_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1907:114
    .z     (_col_5_n_tmp_3_z)
  );
  SHR_14 col_5_n_val_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1624:87
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_tmp_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1623:105
    .z     (_col_5_n_val_3_z)
  );
  CLIP col_5_n_clp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1625:87
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_val_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1624:87
    .z     (n_out_3_5_x)
  );
  SUB col_5_n_tmp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1626:105
    .clock (clock),
    .reset (reset),
    .x     (_col_5_d_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1599:100
    .y     (_delay_INT16_57_1888_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1906:114
    .z     (_col_5_n_tmp_4_z)
  );
  SHR_14 col_5_n_val_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1627:87
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_tmp_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1626:105
    .z     (_col_5_n_val_4_z)
  );
  CLIP col_5_n_clp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1628:87
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_val_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1627:87
    .z     (n_out_4_5_x)
  );
  SUB col_5_n_tmp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1629:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_288_1887_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1905:118
    .y     (_col_5_d_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1613:100
    .z     (_col_5_n_tmp_5_z)
  );
  SHR_14 col_5_n_val_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1630:87
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_tmp_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1629:105
    .z     (_col_5_n_val_5_z)
  );
  CLIP col_5_n_clp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1631:87
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_val_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1630:87
    .z     (n_out_5_5_x)
  );
  SUB col_5_n_tmp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1632:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_180_1886_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1904:118
    .y     (_col_5_d_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1608:100
    .z     (_col_5_n_tmp_6_z)
  );
  SHR_14 col_5_n_val_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1633:87
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_tmp_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1632:105
    .z     (_col_5_n_val_6_z)
  );
  CLIP col_5_n_clp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1634:87
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_val_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1633:87
    .z     (n_out_6_5_x)
  );
  SUB col_5_n_tmp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1635:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_80_2258_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2276:114
    .y     (_col_5_d_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1589:100
    .z     (_col_5_n_tmp_7_z)
  );
  SHR_14 col_5_n_val_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1636:87
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_tmp_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1635:105
    .z     (_col_5_n_val_7_z)
  );
  CLIP col_5_n_clp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1637:87
    .clock (clock),
    .reset (reset),
    .x     (_col_5_n_val_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1636:87
    .z     (n_out_7_5_x)
  );
  C4 col_6_n_c4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1638:70
    .clock (clock),
    .reset (reset),
    .value (_col_6_n_c4_0_value)
  );
  C4 col_6_n_c4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1639:70
    .clock (clock),
    .reset (reset),
    .value (_col_6_n_c4_1_value)
  );
  C4 col_6_n_c4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1640:70
    .clock (clock),
    .reset (reset),
    .value (_col_6_n_c4_2_value)
  );
  C128 col_6_n_c128_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1641:76
    .clock (clock),
    .reset (reset),
    .value (_col_6_n_c128_0_value)
  );
  C128 col_6_n_c128_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1642:76
    .clock (clock),
    .reset (reset),
    .value (_col_6_n_c128_1_value)
  );
  C181 col_6_n_c181_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1643:76
    .clock (clock),
    .reset (reset),
    .value (_col_6_n_c181_0_value)
  );
  C181 col_6_n_c181_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1644:76
    .clock (clock),
    .reset (reset),
    .value (_col_6_n_c181_1_value)
  );
  C8192 col_6_n_c8192 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1645:73
    .clock (clock),
    .reset (reset),
    .value (_col_6_n_c8192_value)
  );
  W7 col_6_n_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1646:64
    .clock (clock),
    .reset (reset),
    .value (_col_6_n_w7_value)
  );
  W1_sub_W7 col_6_n_w1_sub_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1647:85
    .clock (clock),
    .reset (reset),
    .value (_col_6_n_w1_sub_w7_value)
  );
  W1_add_W7 col_6_n_w1_add_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1648:85
    .clock (clock),
    .reset (reset),
    .value (_col_6_n_w1_add_w7_value)
  );
  W3 col_6_n_w3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1649:64
    .clock (clock),
    .reset (reset),
    .value (_col_6_n_w3_value)
  );
  W3_sub_W5 col_6_n_w3_sub_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1650:85
    .clock (clock),
    .reset (reset),
    .value (_col_6_n_w3_sub_w5_value)
  );
  W3_add_W5 col_6_n_w3_add_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1651:85
    .clock (clock),
    .reset (reset),
    .value (_col_6_n_w3_add_w5_value)
  );
  W6 col_6_n_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1652:64
    .clock (clock),
    .reset (reset),
    .value (_col_6_n_w6_value)
  );
  W2_sub_W6 col_6_n_w2_sub_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1653:85
    .clock (clock),
    .reset (reset),
    .value (_col_6_n_w2_sub_w6_value)
  );
  W2_add_W6 col_6_n_w2_add_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1654:85
    .clock (clock),
    .reset (reset),
    .value (_col_6_n_w2_add_w6_value)
  );
  SHL_8 col_6_n_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1655:83
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_shr_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:633:87
    .z     (_col_6_n_x1_0_z)
  );
  SHL_8 col_6_n_t0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1656:83
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_shr_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:241:87
    .z     (_col_6_n_t0_0_z)
  );
  ADD col_6_n_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1657:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_t0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1656:83
    .y     (_col_6_n_c8192_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1645:73
    .z     (_col_6_n_x0_0_z)
  );
  dup_2 col_6_d_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1658:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1657:100
    .y     (_col_6_d_x0_0_y),
    .z     (_col_6_d_x0_0_z)
  );
  dup_2 col_6_d_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1659:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1655:83
    .y     (_col_6_d_x1_0_y),
    .z     (_col_6_d_x1_0_z)
  );
  dup_2 col_6_d_x2_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1660:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_shr_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:829:87
    .y     (_col_6_d_x2_0_y),
    .z     (_col_6_d_x2_0_z)
  );
  dup_2 col_6_d_x3_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1661:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_shr_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:437:87
    .y     (_col_6_d_x3_0_y),
    .z     (_col_6_d_x3_0_z)
  );
  dup_2 col_6_d_x4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1662:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_shr_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:339:87
    .y     (_col_6_d_x4_0_y),
    .z     (_col_6_d_x4_0_z)
  );
  dup_2 col_6_d_x5_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1663:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_shr_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:927:87
    .y     (_col_6_d_x5_0_y),
    .z     (_col_6_d_x5_0_z)
  );
  dup_2 col_6_d_x6_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1664:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_shr_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:731:87
    .y     (_col_6_d_x6_0_y),
    .z     (_col_6_d_x6_0_z)
  );
  dup_2 col_6_d_x7_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1665:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_shr_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:535:87
    .y     (_col_6_d_x7_0_y),
    .z     (_col_6_d_x7_0_z)
  );
  ADD col_6_n_u8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1666:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_11_1885_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1903:114
    .y     (_col_6_d_x5_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1663:100
    .z     (_col_6_n_u8_0_z)
  );
  MUL col_6_n_v8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1667:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1646:64
    .y     (_col_6_n_u8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1666:100
    .z     (_col_6_n_v8_0_z)
  );
  ADD col_6_n_x8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1668:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_v8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1667:100
    .y     (_col_6_n_c4_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1638:70
    .z     (_col_6_n_x8_0_z)
  );
  dup_2 col_6_d_x8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1669:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1668:100
    .y     (_col_6_d_x8_0_y),
    .z     (_col_6_d_x8_0_z)
  );
  MUL col_6_n_u4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1670:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_w1_sub_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1647:85
    .y     (_col_6_d_x4_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1662:100
    .z     (_col_6_n_u4_1_z)
  );
  ADD col_6_n_v4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1671:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_d_x8_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1669:100
    .y     (_delay_INT16_55_1884_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1902:114
    .z     (_col_6_n_v4_1_z)
  );
  SHR_3 col_6_n_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1672:83
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_v4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1671:100
    .z     (_col_6_n_x4_1_z)
  );
  dup_2 col_6_d_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1673:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1672:83
    .y     (_col_6_d_x4_1_y),
    .z     (_col_6_d_x4_1_z)
  );
  MUL col_6_n_u5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1674:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_w1_add_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1648:85
    .y     (_col_6_d_x5_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1663:100
    .z     (_col_6_n_u5_1_z)
  );
  SUB col_6_n_v5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1675:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_d_x8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1669:100
    .y     (_delay_INT16_75_1883_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1901:114
    .z     (_col_6_n_v5_1_z)
  );
  SHR_3 col_6_n_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1676:83
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_v5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1675:100
    .z     (_col_6_n_x5_1_z)
  );
  dup_2 col_6_d_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1677:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1676:83
    .y     (_col_6_d_x5_1_y),
    .z     (_col_6_d_x5_1_z)
  );
  ADD col_6_n_u8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1678:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_d_x6_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1664:100
    .y     (_delay_INT16_1_1948_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1966:110
    .z     (_col_6_n_u8_1_z)
  );
  MUL col_6_n_v8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1679:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_w3_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1649:64
    .y     (_col_6_n_u8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1678:100
    .z     (_col_6_n_v8_1_z)
  );
  ADD col_6_n_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1680:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_v8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1679:100
    .y     (_col_6_n_c4_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1639:70
    .z     (_col_6_n_x8_1_z)
  );
  dup_2 col_6_d_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1681:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1680:100
    .y     (_col_6_d_x8_1_y),
    .z     (_col_6_d_x8_1_z)
  );
  MUL col_6_n_u6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1682:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_w3_sub_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1650:85
    .y     (_col_6_d_x6_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1664:100
    .z     (_col_6_n_u6_1_z)
  );
  SUB col_6_n_v6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1683:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_d_x8_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1681:100
    .y     (_delay_INT16_114_2216_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2234:118
    .z     (_col_6_n_v6_1_z)
  );
  SHR_3 col_6_n_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1684:83
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_v6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1683:100
    .z     (_col_6_n_x6_1_z)
  );
  dup_2 col_6_d_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1685:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1684:83
    .y     (_col_6_d_x6_1_y),
    .z     (_col_6_d_x6_1_z)
  );
  MUL col_6_n_u7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1686:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_w3_add_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1651:85
    .y     (_col_6_d_x7_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1665:100
    .z     (_col_6_n_u7_1_z)
  );
  SUB col_6_n_v7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1687:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_d_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1681:100
    .y     (_delay_INT16_57_2144_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2162:114
    .z     (_col_6_n_v7_1_z)
  );
  SHR_3 col_6_n_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1688:83
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_v7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1687:100
    .z     (_col_6_n_x7_1_z)
  );
  dup_2 col_6_d_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1689:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1688:83
    .y     (_col_6_d_x7_1_y),
    .z     (_col_6_d_x7_1_z)
  );
  ADD col_6_n_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1690:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_d_x0_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1658:100
    .y     (_delay_INT16_5_1882_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1900:110
    .z     (_col_6_n_x8_2_z)
  );
  dup_2 col_6_d_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1691:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1690:100
    .y     (_col_6_d_x8_2_y),
    .z     (_col_6_d_x8_2_z)
  );
  SUB col_6_n_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1692:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_d_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1658:100
    .y     (_delay_INT16_5_2018_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2036:110
    .z     (_col_6_n_x0_1_z)
  );
  dup_2 col_6_d_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1693:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1692:100
    .y     (_col_6_d_x0_1_y),
    .z     (_col_6_d_x0_1_z)
  );
  ADD col_6_n_u1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1694:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_d_x3_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1661:100
    .y     (_delay_INT16_12_1881_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1899:114
    .z     (_col_6_n_u1_1_z)
  );
  MUL col_6_n_v1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1695:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1652:64
    .y     (_col_6_n_u1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1694:100
    .z     (_col_6_n_v1_1_z)
  );
  ADD col_6_n_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1696:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_v1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1695:100
    .y     (_col_6_n_c4_2_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1640:70
    .z     (_col_6_n_x1_1_z)
  );
  dup_2 col_6_d_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1697:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1696:100
    .y     (_col_6_d_x1_1_y),
    .z     (_col_6_d_x1_1_z)
  );
  MUL col_6_n_u2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1698:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_w2_add_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1654:85
    .y     (_col_6_d_x2_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1660:100
    .z     (_col_6_n_u2_1_z)
  );
  SUB col_6_n_v2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1699:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_d_x1_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1697:100
    .y     (_delay_INT16_115_1880_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1898:118
    .z     (_col_6_n_v2_1_z)
  );
  SHR_3 col_6_n_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1700:83
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_v2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1699:100
    .z     (_col_6_n_x2_1_z)
  );
  dup_2 col_6_d_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1701:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1700:83
    .y     (_col_6_d_x2_1_y),
    .z     (_col_6_d_x2_1_z)
  );
  MUL col_6_n_u3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1702:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_w2_sub_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1653:85
    .y     (_col_6_d_x3_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1661:100
    .z     (_col_6_n_u3_1_z)
  );
  ADD col_6_n_v3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1703:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_d_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1697:100
    .y     (_delay_INT16_23_2320_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2338:114
    .z     (_col_6_n_v3_1_z)
  );
  SHR_3 col_6_n_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1704:83
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_v3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1703:100
    .z     (_col_6_n_x3_1_z)
  );
  dup_2 col_6_d_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1705:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1704:83
    .y     (_col_6_d_x3_1_y),
    .z     (_col_6_d_x3_1_z)
  );
  ADD col_6_n_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1706:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_81_2008_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2026:114
    .y     (_col_6_d_x6_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1685:100
    .z     (_col_6_n_x1_2_z)
  );
  dup_2 col_6_d_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1707:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1706:100
    .y     (_col_6_d_x1_2_y),
    .z     (_col_6_d_x1_2_z)
  );
  SUB col_6_n_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1708:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_81_1879_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1897:114
    .y     (_col_6_d_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1685:100
    .z     (_col_6_n_x4_2_z)
  );
  dup_2 col_6_d_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1709:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1708:100
    .y     (_col_6_d_x4_2_y),
    .z     (_col_6_d_x4_2_z)
  );
  ADD col_6_n_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1710:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_d_x5_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1677:100
    .y     (_delay_INT16_83_1878_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1896:114
    .z     (_col_6_n_x6_2_z)
  );
  dup_2 col_6_d_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1711:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1710:100
    .y     (_col_6_d_x6_2_y),
    .z     (_col_6_d_x6_2_z)
  );
  SUB col_6_n_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1712:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_d_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1677:100
    .y     (_delay_INT16_83_2248_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2266:114
    .z     (_col_6_n_x5_2_z)
  );
  dup_2 col_6_d_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1713:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1712:100
    .y     (_col_6_d_x5_2_y),
    .z     (_col_6_d_x5_2_z)
  );
  ADD col_6_n_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1714:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_2_1877_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1895:110
    .y     (_col_6_d_x3_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1705:100
    .z     (_col_6_n_x7_2_z)
  );
  dup_2 col_6_d_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1715:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1714:100
    .y     (_col_6_d_x7_2_y),
    .z     (_col_6_d_x7_2_z)
  );
  SUB col_6_n_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1716:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_2_1960_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1978:110
    .y     (_col_6_d_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1705:100
    .z     (_col_6_n_x8_3_z)
  );
  dup_2 col_6_d_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1717:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1716:100
    .y     (_col_6_d_x8_3_y),
    .z     (_col_6_d_x8_3_z)
  );
  ADD col_6_n_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1718:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_d_x0_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1693:100
    .y     (_delay_INT16_128_1971_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1989:118
    .z     (_col_6_n_x3_2_z)
  );
  dup_2 col_6_d_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1719:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1718:100
    .y     (_col_6_d_x3_2_y),
    .z     (_col_6_d_x3_2_z)
  );
  SUB col_6_n_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1720:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_d_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1693:100
    .y     (_delay_INT16_128_1876_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1894:118
    .z     (_col_6_n_x0_2_z)
  );
  dup_2 col_6_d_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1721:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1720:100
    .y     (_col_6_d_x0_2_y),
    .z     (_col_6_d_x0_2_z)
  );
  ADD col_6_n_u2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1722:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_14_2309_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2327:114
    .y     (_col_6_d_x5_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1713:100
    .z     (_col_6_n_u2_2_z)
  );
  MUL col_6_n_v2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1723:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_c181_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1643:76
    .y     (_col_6_n_u2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1722:100
    .z     (_col_6_n_v2_2_z)
  );
  ADD col_6_n_w2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1724:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_v2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1723:100
    .y     (_col_6_n_c128_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1641:76
    .z     (_col_6_n_w2_2_z)
  );
  SHR_8 col_6_n_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1725:83
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_w2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1724:100
    .z     (_col_6_n_x2_2_z)
  );
  dup_2 col_6_d_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1726:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1725:83
    .y     (_col_6_d_x2_2_y),
    .z     (_col_6_d_x2_2_z)
  );
  SUB col_6_n_u4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1727:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_14_2254_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2272:114
    .y     (_col_6_d_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1713:100
    .z     (_col_6_n_u4_3_z)
  );
  MUL col_6_n_v4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1728:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_c181_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1644:76
    .y     (_col_6_n_u4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1727:100
    .z     (_col_6_n_v4_3_z)
  );
  ADD col_6_n_w4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1729:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_v4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1728:100
    .y     (_col_6_n_c128_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1642:76
    .z     (_col_6_n_w4_3_z)
  );
  SHR_8 col_6_n_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1730:83
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_w4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1729:100
    .z     (_col_6_n_x4_3_z)
  );
  dup_2 col_6_d_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1731:100
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1730:83
    .y     (_col_6_d_x4_3_y),
    .z     (_col_6_d_x4_3_z)
  );
  ADD col_6_n_tmp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1732:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_16_2003_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2021:114
    .y     (_col_6_d_x1_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1707:100
    .z     (_col_6_n_tmp_0_z)
  );
  SHR_14 col_6_n_val_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1733:87
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_tmp_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1732:105
    .z     (_col_6_n_val_0_z)
  );
  CLIP col_6_n_clp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1734:87
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_val_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1733:87
    .z     (n_out_0_6_x)
  );
  ADD col_6_n_tmp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1735:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_106_2054_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2072:118
    .y     (_col_6_d_x2_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1726:100
    .z     (_col_6_n_tmp_1_z)
  );
  SHR_14 col_6_n_val_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1736:87
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_tmp_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1735:105
    .z     (_col_6_n_val_1_z)
  );
  CLIP col_6_n_clp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1737:87
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_val_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1736:87
    .z     (n_out_1_6_x)
  );
  ADD col_6_n_tmp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1738:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_126_1949_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1967:118
    .y     (_col_6_d_x4_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1731:100
    .z     (_col_6_n_tmp_2_z)
  );
  SHR_14 col_6_n_val_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1739:87
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_tmp_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1738:105
    .z     (_col_6_n_val_2_z)
  );
  CLIP col_6_n_clp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1740:87
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_val_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1739:87
    .z     (n_out_2_6_x)
  );
  ADD col_6_n_tmp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1741:105
    .clock (clock),
    .reset (reset),
    .x     (_col_6_d_x8_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1717:100
    .y     (_delay_INT16_29_1875_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1893:114
    .z     (_col_6_n_tmp_3_z)
  );
  SHR_14 col_6_n_val_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1742:87
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_tmp_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1741:105
    .z     (_col_6_n_val_3_z)
  );
  CLIP col_6_n_clp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1743:87
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_val_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1742:87
    .z     (n_out_3_6_x)
  );
  SUB col_6_n_tmp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1744:105
    .clock (clock),
    .reset (reset),
    .x     (_col_6_d_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1717:100
    .y     (_delay_INT16_29_1874_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1892:114
    .z     (_col_6_n_tmp_4_z)
  );
  SHR_14 col_6_n_val_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1745:87
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_tmp_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1744:105
    .z     (_col_6_n_val_4_z)
  );
  CLIP col_6_n_clp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1746:87
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_val_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1745:87
    .z     (n_out_4_6_x)
  );
  SUB col_6_n_tmp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1747:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_126_1873_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1891:118
    .y     (_col_6_d_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1731:100
    .z     (_col_6_n_tmp_5_z)
  );
  SHR_14 col_6_n_val_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1748:87
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_tmp_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1747:105
    .z     (_col_6_n_val_5_z)
  );
  CLIP col_6_n_clp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1749:87
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_val_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1748:87
    .z     (n_out_5_6_x)
  );
  SUB col_6_n_tmp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1750:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_106_1872_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1890:118
    .y     (_col_6_d_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1726:100
    .z     (_col_6_n_tmp_6_z)
  );
  SHR_14 col_6_n_val_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1751:87
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_tmp_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1750:105
    .z     (_col_6_n_val_6_z)
  );
  CLIP col_6_n_clp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1752:87
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_val_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1751:87
    .z     (n_out_6_6_x)
  );
  SUB col_6_n_tmp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1753:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_16_2173_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2191:114
    .y     (_col_6_d_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1707:100
    .z     (_col_6_n_tmp_7_z)
  );
  SHR_14 col_6_n_val_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1754:87
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_tmp_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1753:105
    .z     (_col_6_n_val_7_z)
  );
  CLIP col_6_n_clp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1755:87
    .clock (clock),
    .reset (reset),
    .x     (_col_6_n_val_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1754:87
    .z     (n_out_7_6_x)
  );
  C4 col_7_n_c4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1756:70
    .clock (clock),
    .reset (reset),
    .value (_col_7_n_c4_0_value)
  );
  C4 col_7_n_c4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1757:70
    .clock (clock),
    .reset (reset),
    .value (_col_7_n_c4_1_value)
  );
  C4 col_7_n_c4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1758:70
    .clock (clock),
    .reset (reset),
    .value (_col_7_n_c4_2_value)
  );
  C128 col_7_n_c128_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1759:76
    .clock (clock),
    .reset (reset),
    .value (_col_7_n_c128_0_value)
  );
  C128 col_7_n_c128_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1760:76
    .clock (clock),
    .reset (reset),
    .value (_col_7_n_c128_1_value)
  );
  C181 col_7_n_c181_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1761:76
    .clock (clock),
    .reset (reset),
    .value (_col_7_n_c181_0_value)
  );
  C181 col_7_n_c181_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1762:76
    .clock (clock),
    .reset (reset),
    .value (_col_7_n_c181_1_value)
  );
  C8192 col_7_n_c8192 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1763:73
    .clock (clock),
    .reset (reset),
    .value (_col_7_n_c8192_value)
  );
  W7 col_7_n_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1764:64
    .clock (clock),
    .reset (reset),
    .value (_col_7_n_w7_value)
  );
  W1_sub_W7 col_7_n_w1_sub_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1765:85
    .clock (clock),
    .reset (reset),
    .value (_col_7_n_w1_sub_w7_value)
  );
  W1_add_W7 col_7_n_w1_add_w7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1766:85
    .clock (clock),
    .reset (reset),
    .value (_col_7_n_w1_add_w7_value)
  );
  W3 col_7_n_w3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1767:64
    .clock (clock),
    .reset (reset),
    .value (_col_7_n_w3_value)
  );
  W3_sub_W5 col_7_n_w3_sub_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1768:85
    .clock (clock),
    .reset (reset),
    .value (_col_7_n_w3_sub_w5_value)
  );
  W3_add_W5 col_7_n_w3_add_w5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1769:85
    .clock (clock),
    .reset (reset),
    .value (_col_7_n_w3_add_w5_value)
  );
  W6 col_7_n_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1770:64
    .clock (clock),
    .reset (reset),
    .value (_col_7_n_w6_value)
  );
  W2_sub_W6 col_7_n_w2_sub_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1771:85
    .clock (clock),
    .reset (reset),
    .value (_col_7_n_w2_sub_w6_value)
  );
  W2_add_W6 col_7_n_w2_add_w6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1772:85
    .clock (clock),
    .reset (reset),
    .value (_col_7_n_w2_add_w6_value)
  );
  SHL_8 col_7_n_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1773:83
    .clock (clock),
    .reset (reset),
    .x     (_row_4_n_shr_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:635:87
    .z     (_col_7_n_x1_0_z)
  );
  SHL_8 col_7_n_t0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1774:83
    .clock (clock),
    .reset (reset),
    .x     (_row_0_n_shr_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:243:87
    .z     (_col_7_n_t0_0_z)
  );
  ADD col_7_n_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1775:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_t0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1774:83
    .y     (_col_7_n_c8192_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1763:73
    .z     (_col_7_n_x0_0_z)
  );
  dup_2 col_7_d_x0_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1776:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1775:100
    .y     (_col_7_d_x0_0_y),
    .z     (_col_7_d_x0_0_z)
  );
  dup_2 col_7_d_x1_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1777:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1773:83
    .y     (_col_7_d_x1_0_y),
    .z     (_col_7_d_x1_0_z)
  );
  dup_2 col_7_d_x2_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1778:100
    .clock (clock),
    .reset (reset),
    .x     (_row_6_n_shr_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:831:87
    .y     (_col_7_d_x2_0_y),
    .z     (_col_7_d_x2_0_z)
  );
  dup_2 col_7_d_x3_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1779:100
    .clock (clock),
    .reset (reset),
    .x     (_row_2_n_shr_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:439:87
    .y     (_col_7_d_x3_0_y),
    .z     (_col_7_d_x3_0_z)
  );
  dup_2 col_7_d_x4_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1780:100
    .clock (clock),
    .reset (reset),
    .x     (_row_1_n_shr_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:341:87
    .y     (_col_7_d_x4_0_y),
    .z     (_col_7_d_x4_0_z)
  );
  dup_2 col_7_d_x5_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1781:100
    .clock (clock),
    .reset (reset),
    .x     (_row_7_n_shr_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:929:87
    .y     (_col_7_d_x5_0_y),
    .z     (_col_7_d_x5_0_z)
  );
  dup_2 col_7_d_x6_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1782:100
    .clock (clock),
    .reset (reset),
    .x     (_row_5_n_shr_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:733:87
    .y     (_col_7_d_x6_0_y),
    .z     (_col_7_d_x6_0_z)
  );
  dup_2 col_7_d_x7_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1783:100
    .clock (clock),
    .reset (reset),
    .x     (_row_3_n_shr_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:537:87
    .y     (_col_7_d_x7_0_y),
    .z     (_col_7_d_x7_0_z)
  );
  ADD col_7_n_u8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1784:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_96_1871_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1889:114
    .y     (_col_7_d_x5_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1781:100
    .z     (_col_7_n_u8_0_z)
  );
  MUL col_7_n_v8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1785:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1764:64
    .y     (_col_7_n_u8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1784:100
    .z     (_col_7_n_v8_0_z)
  );
  ADD col_7_n_x8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1786:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_v8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1785:100
    .y     (_col_7_n_c4_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1756:70
    .z     (_col_7_n_x8_0_z)
  );
  dup_2 col_7_d_x8_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1787:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1786:100
    .y     (_col_7_d_x8_0_y),
    .z     (_col_7_d_x8_0_z)
  );
  MUL col_7_n_u4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1788:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_w1_sub_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1765:85
    .y     (_col_7_d_x4_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1780:100
    .z     (_col_7_n_u4_1_z)
  );
  ADD col_7_n_v4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1789:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_d_x8_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1787:100
    .y     (_delay_INT16_245_2286_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2304:118
    .z     (_col_7_n_v4_1_z)
  );
  SHR_3 col_7_n_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1790:83
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_v4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1789:100
    .z     (_col_7_n_x4_1_z)
  );
  dup_2 col_7_d_x4_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1791:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1790:83
    .y     (_col_7_d_x4_1_y),
    .z     (_col_7_d_x4_1_z)
  );
  MUL col_7_n_u5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1792:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_w1_add_w7_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1766:85
    .y     (_col_7_d_x5_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1781:100
    .z     (_col_7_n_u5_1_z)
  );
  SUB col_7_n_v5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1793:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_d_x8_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1787:100
    .y     (_delay_INT16_136_1870_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1888:118
    .z     (_col_7_n_v5_1_z)
  );
  SHR_3 col_7_n_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1794:83
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_v5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1793:100
    .z     (_col_7_n_x5_1_z)
  );
  dup_2 col_7_d_x5_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1795:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1794:83
    .y     (_col_7_d_x5_1_y),
    .z     (_col_7_d_x5_1_z)
  );
  ADD col_7_n_u8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1796:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_d_x6_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1782:100
    .y     (_delay_INT16_78_1869_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1887:114
    .z     (_col_7_n_u8_1_z)
  );
  MUL col_7_n_v8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1797:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_w3_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1767:64
    .y     (_col_7_n_u8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1796:100
    .z     (_col_7_n_v8_1_z)
  );
  ADD col_7_n_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1798:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_v8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1797:100
    .y     (_col_7_n_c4_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1757:70
    .z     (_col_7_n_x8_1_z)
  );
  dup_2 col_7_d_x8_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1799:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1798:100
    .y     (_col_7_d_x8_1_y),
    .z     (_col_7_d_x8_1_z)
  );
  MUL col_7_n_u6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1800:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_w3_sub_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1768:85
    .y     (_col_7_d_x6_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1782:100
    .z     (_col_7_n_u6_1_z)
  );
  SUB col_7_n_v6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1801:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_d_x8_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1799:100
    .y     (_delay_INT16_129_1868_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1886:118
    .z     (_col_7_n_v6_1_z)
  );
  SHR_3 col_7_n_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1802:83
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_v6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1801:100
    .z     (_col_7_n_x6_1_z)
  );
  dup_2 col_7_d_x6_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1803:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1802:83
    .y     (_col_7_d_x6_1_y),
    .z     (_col_7_d_x6_1_z)
  );
  MUL col_7_n_u7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1804:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_w3_add_w5_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1769:85
    .y     (_col_7_d_x7_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1783:100
    .z     (_col_7_n_u7_1_z)
  );
  SUB col_7_n_v7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1805:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_d_x8_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1799:100
    .y     (_delay_INT16_225_2265_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2283:118
    .z     (_col_7_n_v7_1_z)
  );
  SHR_3 col_7_n_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1806:83
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_v7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1805:100
    .z     (_col_7_n_x7_1_z)
  );
  dup_2 col_7_d_x7_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1807:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1806:83
    .y     (_col_7_d_x7_1_y),
    .z     (_col_7_d_x7_1_z)
  );
  ADD col_7_n_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1808:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_68_2112_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2130:114
    .y     (_col_7_d_x1_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1777:100
    .z     (_col_7_n_x8_2_z)
  );
  dup_2 col_7_d_x8_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1809:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1808:100
    .y     (_col_7_d_x8_2_y),
    .z     (_col_7_d_x8_2_z)
  );
  SUB col_7_n_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1810:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_68_2022_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2040:114
    .y     (_col_7_d_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1777:100
    .z     (_col_7_n_x0_1_z)
  );
  dup_2 col_7_d_x0_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1811:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1810:100
    .y     (_col_7_d_x0_1_y),
    .z     (_col_7_d_x0_1_z)
  );
  ADD col_7_n_u1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1812:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_86_1867_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1885:114
    .y     (_col_7_d_x2_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1778:100
    .z     (_col_7_n_u1_1_z)
  );
  MUL col_7_n_v1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1813:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1770:64
    .y     (_col_7_n_u1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1812:100
    .z     (_col_7_n_v1_1_z)
  );
  ADD col_7_n_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1814:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_v1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1813:100
    .y     (_col_7_n_c4_2_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1758:70
    .z     (_col_7_n_x1_1_z)
  );
  dup_2 col_7_d_x1_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1815:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1814:100
    .y     (_col_7_d_x1_1_y),
    .z     (_col_7_d_x1_1_z)
  );
  MUL col_7_n_u2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1816:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_w2_add_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1772:85
    .y     (_col_7_d_x2_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1778:100
    .z     (_col_7_n_u2_1_z)
  );
  SUB col_7_n_v2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1817:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_d_x1_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1815:100
    .y     (_delay_INT16_136_1866_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1884:118
    .z     (_col_7_n_v2_1_z)
  );
  SHR_3 col_7_n_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1818:83
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_v2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1817:100
    .z     (_col_7_n_x2_1_z)
  );
  dup_2 col_7_d_x2_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1819:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1818:83
    .y     (_col_7_d_x2_1_y),
    .z     (_col_7_d_x2_1_z)
  );
  MUL col_7_n_u3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1820:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_w2_sub_w6_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1771:85
    .y     (_col_7_d_x3_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1779:100
    .z     (_col_7_n_u3_1_z)
  );
  ADD col_7_n_v3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1821:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_d_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1815:100
    .y     (_delay_INT16_306_2310_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2328:118
    .z     (_col_7_n_v3_1_z)
  );
  SHR_3 col_7_n_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1822:83
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_v3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1821:100
    .z     (_col_7_n_x3_1_z)
  );
  dup_2 col_7_d_x3_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1823:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1822:83
    .y     (_col_7_d_x3_1_y),
    .z     (_col_7_d_x3_1_z)
  );
  ADD col_7_n_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1824:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_29_2048_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2066:114
    .y     (_col_7_d_x6_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1803:100
    .z     (_col_7_n_x1_2_z)
  );
  dup_2 col_7_d_x1_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1825:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1824:100
    .y     (_col_7_d_x1_2_y),
    .z     (_col_7_d_x1_2_z)
  );
  SUB col_7_n_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1826:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_29_1865_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1883:114
    .y     (_col_7_d_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1803:100
    .z     (_col_7_n_x4_2_z)
  );
  dup_2 col_7_d_x4_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1827:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1826:100
    .y     (_col_7_d_x4_2_y),
    .z     (_col_7_d_x4_2_z)
  );
  ADD col_7_n_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1828:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_d_x5_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1795:100
    .y     (_delay_INT16_1_2080_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2098:110
    .z     (_col_7_n_x6_2_z)
  );
  dup_2 col_7_d_x6_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1829:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1828:100
    .y     (_col_7_d_x6_2_y),
    .z     (_col_7_d_x6_2_z)
  );
  SUB col_7_n_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1830:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_d_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1795:100
    .y     (_delay_INT16_1_1864_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1882:110
    .z     (_col_7_n_x5_2_z)
  );
  dup_2 col_7_d_x5_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1831:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1830:100
    .y     (_col_7_d_x5_2_y),
    .z     (_col_7_d_x5_2_z)
  );
  ADD col_7_n_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1832:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_161_1863_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1881:118
    .y     (_col_7_d_x3_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1823:100
    .z     (_col_7_n_x7_2_z)
  );
  dup_2 col_7_d_x7_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1833:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1832:100
    .y     (_col_7_d_x7_2_y),
    .z     (_col_7_d_x7_2_z)
  );
  SUB col_7_n_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1834:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_161_2189_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2207:118
    .y     (_col_7_d_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1823:100
    .z     (_col_7_n_x8_3_z)
  );
  dup_2 col_7_d_x8_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1835:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1834:100
    .y     (_col_7_d_x8_3_y),
    .z     (_col_7_d_x8_3_z)
  );
  ADD col_7_n_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1836:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_106_1862_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1880:118
    .y     (_col_7_d_x2_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1819:100
    .z     (_col_7_n_x3_2_z)
  );
  dup_2 col_7_d_x3_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1837:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1836:100
    .y     (_col_7_d_x3_2_y),
    .z     (_col_7_d_x3_2_z)
  );
  SUB col_7_n_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1838:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_106_1861_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1879:118
    .y     (_col_7_d_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1819:100
    .z     (_col_7_n_x0_2_z)
  );
  dup_2 col_7_d_x0_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1839:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1838:100
    .y     (_col_7_d_x0_2_y),
    .z     (_col_7_d_x0_2_z)
  );
  ADD col_7_n_u2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1840:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_51_1860_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1878:114
    .y     (_col_7_d_x5_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1831:100
    .z     (_col_7_n_u2_2_z)
  );
  MUL col_7_n_v2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1841:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_c181_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1761:76
    .y     (_col_7_n_u2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1840:100
    .z     (_col_7_n_v2_2_z)
  );
  ADD col_7_n_w2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1842:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_v2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1841:100
    .y     (_col_7_n_c128_0_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1759:76
    .z     (_col_7_n_w2_2_z)
  );
  SHR_8 col_7_n_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1843:83
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_w2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1842:100
    .z     (_col_7_n_x2_2_z)
  );
  dup_2 col_7_d_x2_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1844:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1843:83
    .y     (_col_7_d_x2_2_y),
    .z     (_col_7_d_x2_2_z)
  );
  SUB col_7_n_u4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1845:100
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_51_2156_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2174:114
    .y     (_col_7_d_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1831:100
    .z     (_col_7_n_u4_3_z)
  );
  MUL col_7_n_v4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1846:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_c181_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1762:76
    .y     (_col_7_n_u4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1845:100
    .z     (_col_7_n_v4_3_z)
  );
  ADD col_7_n_w4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1847:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_v4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1846:100
    .y     (_col_7_n_c128_1_value),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1760:76
    .z     (_col_7_n_w4_3_z)
  );
  SHR_8 col_7_n_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1848:83
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_w4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1847:100
    .z     (_col_7_n_x4_3_z)
  );
  dup_2 col_7_d_x4_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1849:100
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1848:83
    .y     (_col_7_d_x4_3_y),
    .z     (_col_7_d_x4_3_z)
  );
  ADD col_7_n_tmp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1850:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_55_2045_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2063:114
    .y     (_col_7_d_x1_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1825:100
    .z     (_col_7_n_tmp_0_z)
  );
  SHR_14 col_7_n_val_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1851:87
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_tmp_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1850:105
    .z     (_col_7_n_val_0_z)
  );
  CLIP col_7_n_clp_0 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1852:87
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_val_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1851:87
    .z     (n_out_0_7_x)
  );
  ADD col_7_n_tmp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1853:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_295_1980_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1998:118
    .y     (_col_7_d_x2_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1844:100
    .z     (_col_7_n_tmp_1_z)
  );
  SHR_14 col_7_n_val_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1854:87
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_tmp_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1853:105
    .z     (_col_7_n_val_1_z)
  );
  CLIP col_7_n_clp_1 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1855:87
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_val_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1854:87
    .z     (n_out_1_7_x)
  );
  ADD col_7_n_tmp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1856:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_397_1978_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1996:118
    .y     (_col_7_d_x4_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1849:100
    .z     (_col_7_n_tmp_2_z)
  );
  SHR_14 col_7_n_val_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1857:87
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_tmp_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1856:105
    .z     (_col_7_n_val_2_z)
  );
  CLIP col_7_n_clp_2 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1858:87
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_val_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1857:87
    .z     (n_out_2_7_x)
  );
  ADD col_7_n_tmp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1859:105
    .clock (clock),
    .reset (reset),
    .x     (_col_7_d_x8_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1835:100
    .y     (_delay_INT16_23_1859_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1877:114
    .z     (_col_7_n_tmp_3_z)
  );
  SHR_14 col_7_n_val_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1860:87
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_tmp_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1859:105
    .z     (_col_7_n_val_3_z)
  );
  CLIP col_7_n_clp_3 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1861:87
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_val_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1860:87
    .z     (n_out_3_7_x)
  );
  SUB col_7_n_tmp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1862:105
    .clock (clock),
    .reset (reset),
    .x     (_col_7_d_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1835:100
    .y     (_delay_INT16_23_1858_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1876:114
    .z     (_col_7_n_tmp_4_z)
  );
  SHR_14 col_7_n_val_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1863:87
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_tmp_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1862:105
    .z     (_col_7_n_val_4_z)
  );
  CLIP col_7_n_clp_4 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1864:87
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_val_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1863:87
    .z     (n_out_4_7_x)
  );
  SUB col_7_n_tmp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1865:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_397_1857_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1875:118
    .y     (_col_7_d_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1849:100
    .z     (_col_7_n_tmp_5_z)
  );
  SHR_14 col_7_n_val_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1866:87
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_tmp_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1865:105
    .z     (_col_7_n_val_5_z)
  );
  CLIP col_7_n_clp_5 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1867:87
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_val_5_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1866:87
    .z     (n_out_5_7_x)
  );
  SUB col_7_n_tmp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1868:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_295_1856_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1874:118
    .y     (_col_7_d_x2_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1844:100
    .z     (_col_7_n_tmp_6_z)
  );
  SHR_14 col_7_n_val_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1869:87
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_tmp_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1868:105
    .z     (_col_7_n_val_6_z)
  );
  CLIP col_7_n_clp_6 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1870:87
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_val_6_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1869:87
    .z     (n_out_6_7_x)
  );
  SUB col_7_n_tmp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1871:105
    .clock (clock),
    .reset (reset),
    .x     (_delay_INT16_55_1938_out),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1956:114
    .y     (_col_7_d_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1825:100
    .z     (_col_7_n_tmp_7_z)
  );
  SHR_14 col_7_n_val_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1872:87
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_tmp_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1871:105
    .z     (_col_7_n_val_7_z)
  );
  CLIP col_7_n_clp_7 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1873:87
    .clock (clock),
    .reset (reset),
    .x     (_col_7_n_val_7_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1872:87
    .z     (n_out_7_7_x)
  );
  delay_INT16_295 delay_INT16_295_1856 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1874:118
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1837:100
    .out   (_delay_INT16_295_1856_out)
  );
  delay_INT16_397 delay_INT16_397_1857 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1875:118
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1839:100
    .out   (_delay_INT16_397_1857_out)
  );
  delay_INT16_23 delay_INT16_23_1858 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1876:114
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1829:100
    .out   (_delay_INT16_23_1858_out)
  );
  delay_INT16_23 delay_INT16_23_1859 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1877:114
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x6_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1829:100
    .out   (_delay_INT16_23_1859_out)
  );
  delay_INT16_51 delay_INT16_51_1860 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1878:114
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x4_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1827:100
    .out   (_delay_INT16_51_1860_out)
  );
  delay_INT16_106 delay_INT16_106_1861 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1879:118
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1811:100
    .out   (_delay_INT16_106_1861_out)
  );
  delay_INT16_106 delay_INT16_106_1862 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1880:118
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x0_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1811:100
    .out   (_delay_INT16_106_1862_out)
  );
  delay_INT16_161 delay_INT16_161_1863 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1881:118
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x8_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1809:100
    .out   (_delay_INT16_161_1863_out)
  );
  delay_INT16_1 delay_INT16_1_1864 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1882:110
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1807:100
    .out   (_delay_INT16_1_1864_out)
  );
  delay_INT16_29 delay_INT16_29_1865 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1883:114
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1791:100
    .out   (_delay_INT16_29_1865_out)
  );
  delay_INT16_136 delay_INT16_136_1866 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1884:118
    .clock (clock),
    .reset (reset),
    .in    (_col_7_n_u2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1816:100
    .out   (_delay_INT16_136_1866_out)
  );
  delay_INT16_86 delay_INT16_86_1867 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1885:114
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x3_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1779:100
    .out   (_delay_INT16_86_1867_out)
  );
  delay_INT16_129 delay_INT16_129_1868 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1886:118
    .clock (clock),
    .reset (reset),
    .in    (_col_7_n_u6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1800:100
    .out   (_delay_INT16_129_1868_out)
  );
  delay_INT16_78 delay_INT16_78_1869 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1887:114
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x7_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1783:100
    .out   (_delay_INT16_78_1869_out)
  );
  delay_INT16_136 delay_INT16_136_1870 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1888:118
    .clock (clock),
    .reset (reset),
    .in    (_col_7_n_u5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1792:100
    .out   (_delay_INT16_136_1870_out)
  );
  delay_INT16_96 delay_INT16_96_1871 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1889:114
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x4_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1780:100
    .out   (_delay_INT16_96_1871_out)
  );
  delay_INT16_106 delay_INT16_106_1872 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1890:118
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1719:100
    .out   (_delay_INT16_106_1872_out)
  );
  delay_INT16_126 delay_INT16_126_1873 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1891:118
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1721:100
    .out   (_delay_INT16_126_1873_out)
  );
  delay_INT16_29 delay_INT16_29_1874 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1892:114
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1711:100
    .out   (_delay_INT16_29_1874_out)
  );
  delay_INT16_29 delay_INT16_29_1875 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1893:114
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x6_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1711:100
    .out   (_delay_INT16_29_1875_out)
  );
  delay_INT16_128 delay_INT16_128_1876 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1894:118
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1701:100
    .out   (_delay_INT16_128_1876_out)
  );
  delay_INT16_2 delay_INT16_2_1877 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1895:110
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x8_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1691:100
    .out   (_delay_INT16_2_1877_out)
  );
  delay_INT16_83 delay_INT16_83_1878 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1896:114
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x7_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1689:100
    .out   (_delay_INT16_83_1878_out)
  );
  delay_INT16_81 delay_INT16_81_1879 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1897:114
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1673:100
    .out   (_delay_INT16_81_1879_out)
  );
  delay_INT16_115 delay_INT16_115_1880 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1898:118
    .clock (clock),
    .reset (reset),
    .in    (_col_6_n_u2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1698:100
    .out   (_delay_INT16_115_1880_out)
  );
  delay_INT16_12 delay_INT16_12_1881 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1899:114
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x2_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1660:100
    .out   (_delay_INT16_12_1881_out)
  );
  delay_INT16_5 delay_INT16_5_1882 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1900:110
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x1_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1659:100
    .out   (_delay_INT16_5_1882_out)
  );
  delay_INT16_75 delay_INT16_75_1883 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1901:114
    .clock (clock),
    .reset (reset),
    .in    (_col_6_n_u5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1674:100
    .out   (_delay_INT16_75_1883_out)
  );
  delay_INT16_55 delay_INT16_55_1884 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1902:114
    .clock (clock),
    .reset (reset),
    .in    (_col_6_n_u4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1670:100
    .out   (_delay_INT16_55_1884_out)
  );
  delay_INT16_11 delay_INT16_11_1885 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1903:114
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x4_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1662:100
    .out   (_delay_INT16_11_1885_out)
  );
  delay_INT16_180 delay_INT16_180_1886 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1904:118
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1601:100
    .out   (_delay_INT16_180_1886_out)
  );
  delay_INT16_288 delay_INT16_288_1887 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1905:118
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1603:100
    .out   (_delay_INT16_288_1887_out)
  );
  delay_INT16_57 delay_INT16_57_1888 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1906:114
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1593:100
    .out   (_delay_INT16_57_1888_out)
  );
  delay_INT16_57 delay_INT16_57_1889 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1907:114
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x6_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1593:100
    .out   (_delay_INT16_57_1889_out)
  );
  delay_INT16_186 delay_INT16_186_1890 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1908:118
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1575:100
    .out   (_delay_INT16_186_1890_out)
  );
  delay_INT16_378 delay_INT16_378_1891 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1909:118
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1555:100
    .out   (_delay_INT16_378_1891_out)
  );
  delay_INT16_126 delay_INT16_126_1892 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1910:118
    .clock (clock),
    .reset (reset),
    .in    (_col_5_n_u2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1580:100
    .out   (_delay_INT16_126_1892_out)
  );
  delay_INT16_81 delay_INT16_81_1893 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1911:114
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x3_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1543:100
    .out   (_delay_INT16_81_1893_out)
  );
  delay_INT16_121 delay_INT16_121_1894 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1912:118
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x0_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1540:100
    .out   (_delay_INT16_121_1894_out)
  );
  delay_INT16_130 delay_INT16_130_1895 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1913:118
    .clock (clock),
    .reset (reset),
    .in    (_col_5_n_u7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1568:100
    .out   (_delay_INT16_130_1895_out)
  );
  delay_INT16_230 delay_INT16_230_1896 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1914:118
    .clock (clock),
    .reset (reset),
    .in    (_col_5_n_u6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1564:100
    .out   (_delay_INT16_230_1896_out)
  );
  delay_INT16_14 delay_INT16_14_1897 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1915:114
    .clock (clock),
    .reset (reset),
    .in    (_col_5_n_u5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1556:100
    .out   (_delay_INT16_14_1897_out)
  );
  delay_INT16_6 delay_INT16_6_1898 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1916:110
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x8_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1551:100
    .out   (_delay_INT16_6_1898_out)
  );
  delay_INT16_26 delay_INT16_26_1899 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1917:114
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x5_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1545:100
    .out   (_delay_INT16_26_1899_out)
  );
  delay_INT16_334 delay_INT16_334_1900 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1918:118
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1485:100
    .out   (_delay_INT16_334_1900_out)
  );
  delay_INT16_2 delay_INT16_2_1901 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1919:110
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1481:100
    .out   (_delay_INT16_2_1901_out)
  );
  delay_INT16_334 delay_INT16_334_1902 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1920:118
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x0_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1485:100
    .out   (_delay_INT16_334_1902_out)
  );
  delay_INT16_38 delay_INT16_38_1903 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1921:114
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x1_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1471:100
    .out   (_delay_INT16_38_1903_out)
  );
  delay_INT16_17 delay_INT16_17_1904 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1922:114
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1465:100
    .out   (_delay_INT16_17_1904_out)
  );
  delay_INT16_21 delay_INT16_21_1905 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1923:114
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x8_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1455:100
    .out   (_delay_INT16_21_1905_out)
  );
  delay_INT16_165 delay_INT16_165_1906 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1924:118
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1453:100
    .out   (_delay_INT16_165_1906_out)
  );
  delay_INT16_165 delay_INT16_165_1907 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1925:118
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x7_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1453:100
    .out   (_delay_INT16_165_1907_out)
  );
  delay_INT16_131 delay_INT16_131_1908 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1926:118
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1449:100
    .out   (_delay_INT16_131_1908_out)
  );
  delay_INT16_159 delay_INT16_159_1909 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1927:118
    .clock (clock),
    .reset (reset),
    .in    (_col_4_n_u3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1466:100
    .out   (_delay_INT16_159_1909_out)
  );
  delay_INT16_207 delay_INT16_207_1910 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1928:118
    .clock (clock),
    .reset (reset),
    .in    (_col_4_n_u2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1462:100
    .out   (_delay_INT16_207_1910_out)
  );
  delay_INT16_351 delay_INT16_351_1911 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1929:118
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1365:100
    .out   (_delay_INT16_351_1911_out)
  );
  delay_INT16_222 delay_INT16_222_1912 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1930:118
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1367:100
    .out   (_delay_INT16_222_1912_out)
  );
  delay_INT16_1 delay_INT16_1_1913 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1931:110
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1363:100
    .out   (_delay_INT16_1_1913_out)
  );
  delay_INT16_1 delay_INT16_1_1914 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1932:110
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x8_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1363:100
    .out   (_delay_INT16_1_1914_out)
  );
  delay_INT16_351 delay_INT16_351_1915 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1933:118
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x3_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1365:100
    .out   (_delay_INT16_351_1915_out)
  );
  delay_INT16_99 delay_INT16_99_1916 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1934:114
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x1_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1353:100
    .out   (_delay_INT16_99_1916_out)
  );
  delay_INT16_27 delay_INT16_27_1917 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1935:114
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x2_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1424:100
    .out   (_delay_INT16_27_1917_out)
  );
  delay_INT16_125 delay_INT16_125_1918 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1936:118
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1422:100
    .out   (_delay_INT16_125_1918_out)
  );
  delay_INT16_125 delay_INT16_125_1919 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1937:118
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x0_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1422:100
    .out   (_delay_INT16_125_1919_out)
  );
  delay_INT16_140 delay_INT16_140_1920 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1938:118
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1355:100
    .out   (_delay_INT16_140_1920_out)
  );
  delay_INT16_106 delay_INT16_106_1921 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1939:118
    .clock (clock),
    .reset (reset),
    .in    (_col_4_n_u7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1450:100
    .out   (_delay_INT16_106_1921_out)
  );
  delay_INT16_140 delay_INT16_140_1922 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1940:118
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x4_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1355:100
    .out   (_delay_INT16_140_1922_out)
  );
  delay_INT16_7 delay_INT16_7_1923 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1941:110
    .clock (clock),
    .reset (reset),
    .in    (_col_4_n_u6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1446:100
    .out   (_delay_INT16_7_1923_out)
  );
  delay_INT16_90 delay_INT16_90_1924 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1942:114
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1339:100
    .out   (_delay_INT16_90_1924_out)
  );
  delay_INT16_90 delay_INT16_90_1925 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1943:114
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x0_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1339:100
    .out   (_delay_INT16_90_1925_out)
  );
  delay_INT16_59 delay_INT16_59_1926 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1944:114
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1337:100
    .out   (_delay_INT16_59_1926_out)
  );
  delay_INT16_59 delay_INT16_59_1927 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1945:114
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x8_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1337:100
    .out   (_delay_INT16_59_1927_out)
  );
  delay_INT16_231 delay_INT16_231_1928 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1946:118
    .clock (clock),
    .reset (reset),
    .in    (_col_4_n_u4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1434:100
    .out   (_delay_INT16_231_1928_out)
  );
  delay_INT16_1 delay_INT16_1_1929 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1947:110
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1331:100
    .out   (_delay_INT16_1_1929_out)
  );
  delay_INT16_1 delay_INT16_1_1930 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1948:110
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x6_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1331:100
    .out   (_delay_INT16_1_1930_out)
  );
  delay_INT16_114 delay_INT16_114_1931 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1949:118
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1305:100
    .out   (_delay_INT16_114_1931_out)
  );
  delay_INT16_114 delay_INT16_114_1932 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1950:118
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x1_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1305:100
    .out   (_delay_INT16_114_1932_out)
  );
  delay_INT16_176 delay_INT16_176_1933 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1951:118
    .clock (clock),
    .reset (reset),
    .in    (_col_3_n_u7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1332:100
    .out   (_delay_INT16_176_1933_out)
  );
  delay_INT16_211 delay_INT16_211_1934 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1952:118
    .clock (clock),
    .reset (reset),
    .in    (_col_3_n_u6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1328:100
    .out   (_delay_INT16_211_1934_out)
  );
  delay_INT16_56 delay_INT16_56_1935 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1953:114
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x6_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1310:100
    .out   (_delay_INT16_56_1935_out)
  );
  delay_INT16_178 delay_INT16_178_1936 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1954:118
    .clock (clock),
    .reset (reset),
    .in    (_col_3_n_u5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1320:100
    .out   (_delay_INT16_178_1936_out)
  );
  delay_INT16_65 delay_INT16_65_1937 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1955:114
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x4_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1308:100
    .out   (_delay_INT16_65_1937_out)
  );
  delay_INT16_55 delay_INT16_55_1938 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1956:114
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1833:100
    .out   (_delay_INT16_55_1938_out)
  );
  delay_INT16_122 delay_INT16_122_1939 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1957:118
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1235:100
    .out   (_delay_INT16_122_1939_out)
  );
  delay_INT16_121 delay_INT16_121_1940 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1958:118
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1247:100
    .out   (_delay_INT16_121_1940_out)
  );
  delay_INT16_110 delay_INT16_110_1941 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1959:118
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1249:100
    .out   (_delay_INT16_110_1941_out)
  );
  delay_INT16_145 delay_INT16_145_1942 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1960:118
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x6_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1239:100
    .out   (_delay_INT16_145_1942_out)
  );
  delay_INT16_110 delay_INT16_110_1943 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1961:118
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x0_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1249:100
    .out   (_delay_INT16_110_1943_out)
  );
  delay_INT16_121 delay_INT16_121_1944 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1962:118
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x3_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1247:100
    .out   (_delay_INT16_121_1944_out)
  );
  delay_INT16_122 delay_INT16_122_1945 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1963:118
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x1_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1235:100
    .out   (_delay_INT16_122_1945_out)
  );
  delay_INT16_90 delay_INT16_90_1946 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1964:114
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1241:100
    .out   (_delay_INT16_90_1946_out)
  );
  delay_INT16_378 delay_INT16_378_1947 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1965:118
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x5_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1559:100
    .out   (_delay_INT16_378_1947_out)
  );
  delay_INT16_1 delay_INT16_1_1948 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1966:110
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x7_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1665:100
    .out   (_delay_INT16_1_1948_out)
  );
  delay_INT16_126 delay_INT16_126_1949 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1967:118
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x0_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1721:100
    .out   (_delay_INT16_126_1949_out)
  );
  delay_INT16_66 delay_INT16_66_1950 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1968:114
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x0_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1221:100
    .out   (_delay_INT16_66_1950_out)
  );
  delay_INT16_75 delay_INT16_75_1951 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1969:114
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1233:100
    .out   (_delay_INT16_75_1951_out)
  );
  delay_INT16_64 delay_INT16_64_1952 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1970:114
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1205:100
    .out   (_delay_INT16_64_1952_out)
  );
  delay_INT16_168 delay_INT16_168_1953 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1971:118
    .clock (clock),
    .reset (reset),
    .in    (_col_2_n_u3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1230:100
    .out   (_delay_INT16_168_1953_out)
  );
  delay_INT16_66 delay_INT16_66_1954 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1972:114
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x3_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1189:100
    .out   (_delay_INT16_66_1954_out)
  );
  delay_INT16_213 delay_INT16_213_1955 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1973:118
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x0_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1186:100
    .out   (_delay_INT16_213_1955_out)
  );
  delay_INT16_131 delay_INT16_131_1956 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1974:118
    .clock (clock),
    .reset (reset),
    .in    (_col_2_n_u7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1214:100
    .out   (_delay_INT16_131_1956_out)
  );
  delay_INT16_68 delay_INT16_68_1957 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1975:114
    .clock (clock),
    .reset (reset),
    .in    (_col_2_n_u5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1202:100
    .out   (_delay_INT16_68_1957_out)
  );
  delay_INT16_112 delay_INT16_112_1958 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1976:118
    .clock (clock),
    .reset (reset),
    .in    (_col_2_n_u4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1198:100
    .out   (_delay_INT16_112_1958_out)
  );
  delay_INT16_34 delay_INT16_34_1959 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1977:114
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x4_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1190:100
    .out   (_delay_INT16_34_1959_out)
  );
  delay_INT16_2 delay_INT16_2_1960 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1978:110
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1691:100
    .out   (_delay_INT16_2_1960_out)
  );
  delay_INT16_1 delay_INT16_1_1961 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1979:110
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1117:100
    .out   (_delay_INT16_1_1961_out)
  );
  delay_INT16_190 delay_INT16_190_1962 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1980:118
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1129:100
    .out   (_delay_INT16_190_1962_out)
  );
  delay_INT16_19 delay_INT16_19_1963 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1981:114
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x4_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1141:100
    .out   (_delay_INT16_19_1963_out)
  );
  delay_INT16_73 delay_INT16_73_1964 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1982:114
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x6_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1121:100
    .out   (_delay_INT16_73_1964_out)
  );
  delay_INT16_190 delay_INT16_190_1965 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1983:118
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x3_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1129:100
    .out   (_delay_INT16_190_1965_out)
  );
  delay_INT16_1 delay_INT16_1_1966 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1984:110
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x1_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1117:100
    .out   (_delay_INT16_1_1966_out)
  );
  delay_INT16_17 delay_INT16_17_1967 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1985:114
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x2_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1465:100
    .out   (_delay_INT16_17_1967_out)
  );
  delay_INT16_2 delay_INT16_2_1968 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1986:110
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x4_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1119:100
    .out   (_delay_INT16_2_1968_out)
  );
  delay_INT16_45 delay_INT16_45_1969 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1987:114
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1103:100
    .out   (_delay_INT16_45_1969_out)
  );
  delay_INT16_45 delay_INT16_45_1970 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1988:114
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x0_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1103:100
    .out   (_delay_INT16_45_1970_out)
  );
  delay_INT16_128 delay_INT16_128_1971 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1989:118
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x2_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1701:100
    .out   (_delay_INT16_128_1971_out)
  );
  delay_INT16_27 delay_INT16_27_1972 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1990:114
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1115:100
    .out   (_delay_INT16_27_1972_out)
  );
  delay_INT16_27 delay_INT16_27_1973 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1991:114
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x3_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1115:100
    .out   (_delay_INT16_27_1973_out)
  );
  delay_INT16_10 delay_INT16_10_1974 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1992:114
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1099:100
    .out   (_delay_INT16_10_1974_out)
  );
  delay_INT16_10 delay_INT16_10_1975 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1993:114
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x7_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1099:100
    .out   (_delay_INT16_10_1975_out)
  );
  delay_INT16_64 delay_INT16_64_1976 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1994:114
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1095:100
    .out   (_delay_INT16_64_1976_out)
  );
  delay_INT16_109 delay_INT16_109_1977 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1995:118
    .clock (clock),
    .reset (reset),
    .in    (_col_1_n_u2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1108:100
    .out   (_delay_INT16_109_1977_out)
  );
  delay_INT16_397 delay_INT16_397_1978 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1996:118
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x0_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1839:100
    .out   (_delay_INT16_397_1978_out)
  );
  delay_INT16_131 delay_INT16_131_1979 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1997:118
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1069:100
    .out   (_delay_INT16_131_1979_out)
  );
  delay_INT16_295 delay_INT16_295_1980 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1998:118
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x3_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1837:100
    .out   (_delay_INT16_295_1980_out)
  );
  delay_INT16_131 delay_INT16_131_1981 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1999:118
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x1_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1069:100
    .out   (_delay_INT16_131_1981_out)
  );
  delay_INT16_102 delay_INT16_102_1982 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2000:118
    .clock (clock),
    .reset (reset),
    .in    (_col_1_n_u7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1096:100
    .out   (_delay_INT16_102_1982_out)
  );
  delay_INT16_191 delay_INT16_191_1983 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2001:118
    .clock (clock),
    .reset (reset),
    .in    (_col_1_n_u6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1092:100
    .out   (_delay_INT16_191_1983_out)
  );
  delay_INT16_259 delay_INT16_259_1984 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2002:118
    .clock (clock),
    .reset (reset),
    .in    (_col_1_n_u3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1112:100
    .out   (_delay_INT16_259_1984_out)
  );
  delay_INT16_88 delay_INT16_88_1985 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2003:114
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x6_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1074:100
    .out   (_delay_INT16_88_1985_out)
  );
  delay_INT16_90 delay_INT16_90_1986 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2004:114
    .clock (clock),
    .reset (reset),
    .in    (_col_1_n_u5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1084:100
    .out   (_delay_INT16_90_1986_out)
  );
  delay_INT16_262 delay_INT16_262_1987 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2005:118
    .clock (clock),
    .reset (reset),
    .in    (_col_1_n_u4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1080:100
    .out   (_delay_INT16_262_1987_out)
  );
  delay_INT16_129 delay_INT16_129_1988 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2006:118
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x4_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1072:100
    .out   (_delay_INT16_129_1988_out)
  );
  delay_INT16_213 delay_INT16_213_1989 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2007:118
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1186:100
    .out   (_delay_INT16_213_1989_out)
  );
  delay_INT16_94 delay_INT16_94_1990 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2008:114
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1007:100
    .out   (_delay_INT16_94_1990_out)
  );
  delay_INT16_487 delay_INT16_487_1991 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2009:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1011:100
    .out   (_delay_INT16_487_1991_out)
  );
  delay_INT16_477 delay_INT16_477_1992 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2010:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1013:100
    .out   (_delay_INT16_477_1992_out)
  );
  delay_INT16_34 delay_INT16_34_1993 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2011:114
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x6_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1003:100
    .out   (_delay_INT16_34_1993_out)
  );
  delay_INT16_487 delay_INT16_487_1994 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2012:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x3_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1011:100
    .out   (_delay_INT16_487_1994_out)
  );
  delay_INT16_94 delay_INT16_94_1995 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2013:114
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x7_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1007:100
    .out   (_delay_INT16_94_1995_out)
  );
  delay_INT16_89 delay_INT16_89_1996 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2014:114
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1005:100
    .out   (_delay_INT16_89_1996_out)
  );
  delay_INT16_89 delay_INT16_89_1997 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2015:114
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x5_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1005:100
    .out   (_delay_INT16_89_1997_out)
  );
  delay_INT16_23 delay_INT16_23_1998 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2016:114
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:985:100
    .out   (_delay_INT16_23_1998_out)
  );
  delay_INT16_23 delay_INT16_23_1999 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2017:114
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x0_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:985:100
    .out   (_delay_INT16_23_1999_out)
  );
  delay_INT16_139 delay_INT16_139_2000 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2018:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:983:100
    .out   (_delay_INT16_139_2000_out)
  );
  delay_INT16_139 delay_INT16_139_2001 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2019:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x8_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:983:100
    .out   (_delay_INT16_139_2001_out)
  );
  delay_INT16_94 delay_INT16_94_2002 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2020:114
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:969:100
    .out   (_delay_INT16_94_2002_out)
  );
  delay_INT16_16 delay_INT16_16_2003 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2021:114
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x7_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1715:100
    .out   (_delay_INT16_16_2003_out)
  );
  delay_INT16_94 delay_INT16_94_2004 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2022:114
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x5_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:969:100
    .out   (_delay_INT16_94_2004_out)
  );
  delay_INT16_21 delay_INT16_21_2005 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2023:114
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1455:100
    .out   (_delay_INT16_21_2005_out)
  );
  delay_INT16_212 delay_INT16_212_2006 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2024:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:965:100
    .out   (_delay_INT16_212_2006_out)
  );
  delay_INT16_212 delay_INT16_212_2007 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2025:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x4_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:965:100
    .out   (_delay_INT16_212_2007_out)
  );
  delay_INT16_81 delay_INT16_81_2008 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2026:114
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x4_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1673:100
    .out   (_delay_INT16_81_2008_out)
  );
  delay_INT16_296 delay_INT16_296_2009 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2027:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_n_u3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:994:100
    .out   (_delay_INT16_296_2009_out)
  );
  delay_INT16_90 delay_INT16_90_2010 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2028:114
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x5_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1241:100
    .out   (_delay_INT16_90_2010_out)
  );
  delay_INT16_127 delay_INT16_127_2011 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2029:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_n_u2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:990:100
    .out   (_delay_INT16_127_2011_out)
  );
  delay_INT16_242 delay_INT16_242_2012 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2030:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:950:100
    .out   (_delay_INT16_242_2012_out)
  );
  delay_INT16_338 delay_INT16_338_2013 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2031:118
    .clock (clock),
    .reset (reset),
    .in    (_col_3_n_u2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1344:100
    .out   (_delay_INT16_338_2013_out)
  );
  delay_INT16_242 delay_INT16_242_2014 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2032:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x0_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:950:100
    .out   (_delay_INT16_242_2014_out)
  );
  delay_INT16_145 delay_INT16_145_2015 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2033:118
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1239:100
    .out   (_delay_INT16_145_2015_out)
  );
  delay_INT16_181 delay_INT16_181_2016 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2034:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x6_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:956:100
    .out   (_delay_INT16_181_2016_out)
  );
  delay_INT16_298 delay_INT16_298_2017 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2035:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_n_u5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:966:100
    .out   (_delay_INT16_298_2017_out)
  );
  delay_INT16_5 delay_INT16_5_2018 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2036:110
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1659:100
    .out   (_delay_INT16_5_2018_out)
  );
  delay_INT16_7 delay_INT16_7_2019 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2037:110
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x4_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:954:100
    .out   (_delay_INT16_7_2019_out)
  );
  delay_INT16_64 delay_INT16_64_2020 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2038:114
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x6_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1095:100
    .out   (_delay_INT16_64_2020_out)
  );
  delay_INT16_156 delay_INT16_156_2021 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2039:118
    .clock (clock),
    .reset (reset),
    .in    (_col_2_n_u2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1226:100
    .out   (_delay_INT16_156_2021_out)
  );
  delay_INT16_68 delay_INT16_68_2022 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2040:114
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1776:100
    .out   (_delay_INT16_68_2022_out)
  );
  delay_INT16_45 delay_INT16_45_2023 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2041:114
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:897:100
    .out   (_delay_INT16_45_2023_out)
  );
  delay_INT16_338 delay_INT16_338_2024 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2042:118
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:901:100
    .out   (_delay_INT16_338_2024_out)
  );
  delay_INT16_38 delay_INT16_38_2025 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2043:114
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1471:100
    .out   (_delay_INT16_38_2025_out)
  );
  delay_INT16_255 delay_INT16_255_2026 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2044:118
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:903:100
    .out   (_delay_INT16_255_2026_out)
  );
  delay_INT16_122 delay_INT16_122_2027 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2045:118
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:893:100
    .out   (_delay_INT16_122_2027_out)
  );
  delay_INT16_122 delay_INT16_122_2028 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2046:118
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x6_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:893:100
    .out   (_delay_INT16_122_2028_out)
  );
  delay_INT16_255 delay_INT16_255_2029 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2047:118
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x0_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:903:100
    .out   (_delay_INT16_255_2029_out)
  );
  delay_INT16_338 delay_INT16_338_2030 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2048:118
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x3_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:901:100
    .out   (_delay_INT16_338_2030_out)
  );
  delay_INT16_45 delay_INT16_45_2031 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2049:114
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x7_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:897:100
    .out   (_delay_INT16_45_2031_out)
  );
  delay_INT16_13 delay_INT16_13_2032 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2050:114
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:895:100
    .out   (_delay_INT16_13_2032_out)
  );
  delay_INT16_13 delay_INT16_13_2033 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2051:114
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x5_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:895:100
    .out   (_delay_INT16_13_2033_out)
  );
  delay_INT16_288 delay_INT16_288_2034 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2052:118
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x0_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1603:100
    .out   (_delay_INT16_288_2034_out)
  );
  delay_INT16_19 delay_INT16_19_2035 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2053:114
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x0_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:878:100
    .out   (_delay_INT16_19_2035_out)
  );
  delay_INT16_6 delay_INT16_6_2036 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2054:110
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:887:100
    .out   (_delay_INT16_6_2036_out)
  );
  delay_INT16_35 delay_INT16_35_2037 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2055:114
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:865:100
    .out   (_delay_INT16_35_2037_out)
  );
  delay_INT16_35 delay_INT16_35_2038 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2056:114
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x5_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:865:100
    .out   (_delay_INT16_35_2038_out)
  );
  delay_INT16_33 delay_INT16_33_2039 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2057:114
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x4_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:862:100
    .out   (_delay_INT16_33_2039_out)
  );
  delay_INT16_100 delay_INT16_100_2040 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2058:118
    .clock (clock),
    .reset (reset),
    .in    (_row_7_n_t2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:882:100
    .out   (_delay_INT16_100_2040_out)
  );
  delay_INT16_13 delay_INT16_13_2041 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2059:114
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x2_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:851:100
    .out   (_delay_INT16_13_2041_out)
  );
  delay_INT16_133 delay_INT16_133_2042 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2060:118
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x2_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1306:100
    .out   (_delay_INT16_133_2042_out)
  );
  delay_INT16_121 delay_INT16_121_2043 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2061:118
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x2_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:851:100
    .out   (_delay_INT16_121_2043_out)
  );
  delay_INT16_48 delay_INT16_48_2044 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2062:114
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:849:100
    .out   (_delay_INT16_48_2044_out)
  );
  delay_INT16_55 delay_INT16_55_2045 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2063:114
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x7_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1833:100
    .out   (_delay_INT16_55_2045_out)
  );
  delay_INT16_147 delay_INT16_147_2046 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2064:118
    .clock (clock),
    .reset (reset),
    .in    (_row_7_n_t7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:872:100
    .out   (_delay_INT16_147_2046_out)
  );
  delay_INT16_182 delay_INT16_182_2047 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2065:118
    .clock (clock),
    .reset (reset),
    .in    (_row_7_n_t6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:869:100
    .out   (_delay_INT16_182_2047_out)
  );
  delay_INT16_29 delay_INT16_29_2048 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2066:114
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x4_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1791:100
    .out   (_delay_INT16_29_2048_out)
  );
  delay_INT16_1 delay_INT16_1_2049 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2067:110
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x7_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:856:100
    .out   (_delay_INT16_1_2049_out)
  );
  delay_INT16_111 delay_INT16_111_2050 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2068:118
    .clock (clock),
    .reset (reset),
    .in    (_row_7_n_t5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:863:100
    .out   (_delay_INT16_111_2050_out)
  );
  delay_INT16_187 delay_INT16_187_2051 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2069:118
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x5_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1323:100
    .out   (_delay_INT16_187_2051_out)
  );
  delay_INT16_62 delay_INT16_62_2052 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2070:114
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x3_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1071:100
    .out   (_delay_INT16_62_2052_out)
  );
  delay_INT16_34 delay_INT16_34_2053 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2071:114
    .clock (clock),
    .reset (reset),
    .in    (_row_7_n_t4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:860:100
    .out   (_delay_INT16_34_2053_out)
  );
  delay_INT16_106 delay_INT16_106_2054 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2072:118
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x3_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1719:100
    .out   (_delay_INT16_106_2054_out)
  );
  delay_INT16_19 delay_INT16_19_2055 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2073:114
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x5_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:854:100
    .out   (_delay_INT16_19_2055_out)
  );
  delay_INT16_50 delay_INT16_50_2056 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2074:114
    .clock (clock),
    .reset (reset),
    .in    (_col_2_n_u6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1210:100
    .out   (_delay_INT16_50_2056_out)
  );
  delay_INT16_396 delay_INT16_396_2057 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2075:118
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:803:100
    .out   (_delay_INT16_396_2057_out)
  );
  delay_INT16_2 delay_INT16_2_2058 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2076:110
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x8_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1481:100
    .out   (_delay_INT16_2_2058_out)
  );
  delay_INT16_339 delay_INT16_339_2059 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2077:118
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:805:100
    .out   (_delay_INT16_339_2059_out)
  );
  delay_INT16_142 delay_INT16_142_2060 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2078:118
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x8_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:801:100
    .out   (_delay_INT16_142_2060_out)
  );
  delay_INT16_142 delay_INT16_142_2061 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2079:118
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x8_4_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:801:100
    .out   (_delay_INT16_142_2061_out)
  );
  delay_INT16_396 delay_INT16_396_2062 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2080:118
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x3_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:803:100
    .out   (_delay_INT16_396_2062_out)
  );
  delay_INT16_120 delay_INT16_120_2063 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2081:118
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x7_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:799:100
    .out   (_delay_INT16_120_2063_out)
  );
  delay_INT16_68 delay_INT16_68_2064 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2082:114
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x5_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:797:100
    .out   (_delay_INT16_68_2064_out)
  );
  delay_INT16_14 delay_INT16_14_2065 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2083:114
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:786:100
    .out   (_delay_INT16_14_2065_out)
  );
  delay_INT16_14 delay_INT16_14_2066 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2084:114
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x2_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:786:100
    .out   (_delay_INT16_14_2066_out)
  );
  delay_INT16_15 delay_INT16_15_2067 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2085:114
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:789:100
    .out   (_delay_INT16_15_2067_out)
  );
  delay_INT16_15 delay_INT16_15_2068 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2086:114
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x3_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:789:100
    .out   (_delay_INT16_15_2068_out)
  );
  delay_INT16_17 delay_INT16_17_2069 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2087:114
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:776:100
    .out   (_delay_INT16_17_2069_out)
  );
  delay_INT16_17 delay_INT16_17_2070 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2088:114
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x7_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:776:100
    .out   (_delay_INT16_17_2070_out)
  );
  delay_INT16_24 delay_INT16_24_2071 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2089:114
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:773:100
    .out   (_delay_INT16_24_2071_out)
  );
  delay_INT16_24 delay_INT16_24_2072 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2090:114
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x6_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:773:100
    .out   (_delay_INT16_24_2072_out)
  );
  delay_INT16_99 delay_INT16_99_2073 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2091:114
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1353:100
    .out   (_delay_INT16_99_2073_out)
  );
  delay_INT16_11 delay_INT16_11_2074 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2092:114
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x1_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:783:100
    .out   (_delay_INT16_11_2074_out)
  );
  delay_INT16_17 delay_INT16_17_2075 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2093:114
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x3_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:754:100
    .out   (_delay_INT16_17_2075_out)
  );
  delay_INT16_39 delay_INT16_39_2076 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2094:114
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x1_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:752:100
    .out   (_delay_INT16_39_2076_out)
  );
  delay_INT16_3 delay_INT16_3_2077 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2095:110
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x7_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:758:100
    .out   (_delay_INT16_3_2077_out)
  );
  delay_INT16_173 delay_INT16_173_2078 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2096:118
    .clock (clock),
    .reset (reset),
    .in    (_row_6_n_t5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:765:100
    .out   (_delay_INT16_173_2078_out)
  );
  delay_INT16_47 delay_INT16_47_2079 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2097:114
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x4_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:755:100
    .out   (_delay_INT16_47_2079_out)
  );
  delay_INT16_1 delay_INT16_1_2080 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2098:110
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x7_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1807:100
    .out   (_delay_INT16_1_2080_out)
  );
  delay_INT16_2 delay_INT16_2_2081 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2099:110
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1119:100
    .out   (_delay_INT16_2_2081_out)
  );
  delay_INT16_24 delay_INT16_24_2082 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2100:114
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x5_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1595:100
    .out   (_delay_INT16_24_2082_out)
  );
  delay_INT16_131 delay_INT16_131_2083 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2101:118
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x6_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1449:100
    .out   (_delay_INT16_131_2083_out)
  );
  delay_INT16_134 delay_INT16_134_2084 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2102:118
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:705:100
    .out   (_delay_INT16_134_2084_out)
  );
  delay_INT16_134 delay_INT16_134_2085 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2103:118
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:707:100
    .out   (_delay_INT16_134_2085_out)
  );
  delay_INT16_134 delay_INT16_134_2086 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2104:118
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x0_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:707:100
    .out   (_delay_INT16_134_2086_out)
  );
  delay_INT16_134 delay_INT16_134_2087 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2105:118
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x3_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:705:100
    .out   (_delay_INT16_134_2087_out)
  );
  delay_INT16_142 delay_INT16_142_2088 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2106:118
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x1_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:693:100
    .out   (_delay_INT16_142_2088_out)
  );
  delay_INT16_63 delay_INT16_63_2089 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2107:114
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x4_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:695:100
    .out   (_delay_INT16_63_2089_out)
  );
  delay_INT16_141 delay_INT16_141_2090 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2108:118
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:682:100
    .out   (_delay_INT16_141_2090_out)
  );
  delay_INT16_78 delay_INT16_78_2091 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2109:114
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1201:100
    .out   (_delay_INT16_78_2091_out)
  );
  delay_INT16_115 delay_INT16_115_2092 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2110:118
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x8_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:680:100
    .out   (_delay_INT16_115_2092_out)
  );
  delay_INT16_33 delay_INT16_33_2093 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2111:114
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:862:100
    .out   (_delay_INT16_33_2093_out)
  );
  delay_INT16_61 delay_INT16_61_2094 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2112:114
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:678:100
    .out   (_delay_INT16_61_2094_out)
  );
  delay_INT16_61 delay_INT16_61_2095 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2113:114
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x7_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:678:100
    .out   (_delay_INT16_61_2095_out)
  );
  delay_INT16_5 delay_INT16_5_2096 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2114:110
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:675:100
    .out   (_delay_INT16_5_2096_out)
  );
  delay_INT16_24 delay_INT16_24_2097 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2115:114
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1595:100
    .out   (_delay_INT16_24_2097_out)
  );
  delay_INT16_5 delay_INT16_5_2098 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2116:110
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x6_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:675:100
    .out   (_delay_INT16_5_2098_out)
  );
  delay_INT16_224 delay_INT16_224_2099 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2117:118
    .clock (clock),
    .reset (reset),
    .in    (_row_5_n_t3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:689:100
    .out   (_delay_INT16_224_2099_out)
  );
  delay_INT16_226 delay_INT16_226_2100 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2118:118
    .clock (clock),
    .reset (reset),
    .in    (_row_5_n_t2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:686:100
    .out   (_delay_INT16_226_2100_out)
  );
  delay_INT16_31 delay_INT16_31_2101 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2119:114
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x2_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:655:100
    .out   (_delay_INT16_31_2101_out)
  );
  delay_INT16_8 delay_INT16_8_2102 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2120:110
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:653:100
    .out   (_delay_INT16_8_2102_out)
  );
  delay_INT16_8 delay_INT16_8_2103 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2121:110
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x0_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:653:100
    .out   (_delay_INT16_8_2103_out)
  );
  delay_INT16_87 delay_INT16_87_2104 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2122:114
    .clock (clock),
    .reset (reset),
    .in    (_row_5_n_t7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:676:100
    .out   (_delay_INT16_87_2104_out)
  );
  delay_INT16_43 delay_INT16_43_2105 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2123:114
    .clock (clock),
    .reset (reset),
    .in    (_row_5_n_t6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:673:100
    .out   (_delay_INT16_43_2105_out)
  );
  delay_INT16_10 delay_INT16_10_2106 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2124:114
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x7_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:660:100
    .out   (_delay_INT16_10_2106_out)
  );
  delay_INT16_121 delay_INT16_121_2107 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2125:118
    .clock (clock),
    .reset (reset),
    .in    (_row_5_n_t5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:667:100
    .out   (_delay_INT16_121_2107_out)
  );
  delay_INT16_13 delay_INT16_13_2108 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2126:114
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x5_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:658:100
    .out   (_delay_INT16_13_2108_out)
  );
  delay_INT16_10 delay_INT16_10_2109 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2127:114
    .clock (clock),
    .reset (reset),
    .in    (_row_5_n_t4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:664:100
    .out   (_delay_INT16_10_2109_out)
  );
  delay_INT16_87 delay_INT16_87_2110 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2128:114
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x5_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:658:100
    .out   (_delay_INT16_87_2110_out)
  );
  delay_INT16_73 delay_INT16_73_2111 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2129:114
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1121:100
    .out   (_delay_INT16_73_2111_out)
  );
  delay_INT16_68 delay_INT16_68_2112 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2130:114
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x0_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1776:100
    .out   (_delay_INT16_68_2112_out)
  );
  delay_INT16_83 delay_INT16_83_2113 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2131:114
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:595:100
    .out   (_delay_INT16_83_2113_out)
  );
  delay_INT16_248 delay_INT16_248_2114 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2132:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:607:100
    .out   (_delay_INT16_248_2114_out)
  );
  delay_INT16_222 delay_INT16_222_2115 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2133:118
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x0_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1367:100
    .out   (_delay_INT16_222_2115_out)
  );
  delay_INT16_141 delay_INT16_141_2116 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2134:118
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x0_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:682:100
    .out   (_delay_INT16_141_2116_out)
  );
  delay_INT16_350 delay_INT16_350_2117 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2135:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x0_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:609:100
    .out   (_delay_INT16_350_2117_out)
  );
  delay_INT16_248 delay_INT16_248_2118 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2136:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x3_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:607:100
    .out   (_delay_INT16_248_2118_out)
  );
  delay_INT16_83 delay_INT16_83_2119 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2137:114
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x1_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:595:100
    .out   (_delay_INT16_83_2119_out)
  );
  delay_INT16_114 delay_INT16_114_2120 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2138:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:597:100
    .out   (_delay_INT16_114_2120_out)
  );
  delay_INT16_66 delay_INT16_66_2121 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2139:114
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1221:100
    .out   (_delay_INT16_66_2121_out)
  );
  delay_INT16_114 delay_INT16_114_2122 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2140:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x4_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:597:100
    .out   (_delay_INT16_114_2122_out)
  );
  delay_INT16_370 delay_INT16_370_2123 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2141:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_n_u6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:974:100
    .out   (_delay_INT16_370_2123_out)
  );
  delay_INT16_166 delay_INT16_166_2124 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2142:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:584:100
    .out   (_delay_INT16_166_2124_out)
  );
  delay_INT16_166 delay_INT16_166_2125 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2143:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x0_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:584:100
    .out   (_delay_INT16_166_2125_out)
  );
  delay_INT16_229 delay_INT16_229_2126 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2144:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:582:100
    .out   (_delay_INT16_229_2126_out)
  );
  delay_INT16_117 delay_INT16_117_2127 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2145:118
    .clock (clock),
    .reset (reset),
    .in    (_row_6_n_t7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:774:100
    .out   (_delay_INT16_117_2127_out)
  );
  delay_INT16_229 delay_INT16_229_2128 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2146:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x8_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:582:100
    .out   (_delay_INT16_229_2128_out)
  );
  delay_INT16_95 delay_INT16_95_2129 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2147:114
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:571:100
    .out   (_delay_INT16_95_2129_out)
  );
  delay_INT16_95 delay_INT16_95_2130 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2148:114
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x5_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:571:100
    .out   (_delay_INT16_95_2130_out)
  );
  delay_INT16_79 delay_INT16_79_2131 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2149:114
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:568:100
    .out   (_delay_INT16_79_2131_out)
  );
  delay_INT16_79 delay_INT16_79_2132 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2150:114
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x4_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:568:100
    .out   (_delay_INT16_79_2132_out)
  );
  delay_INT16_68 delay_INT16_68_2133 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2151:114
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x5_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:797:100
    .out   (_delay_INT16_68_2133_out)
  );
  delay_INT16_145 delay_INT16_145_2134 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2152:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_n_t2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:588:100
    .out   (_delay_INT16_145_2134_out)
  );
  delay_INT16_185 delay_INT16_185_2135 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2153:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_n_u7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:978:100
    .out   (_delay_INT16_185_2135_out)
  );
  delay_INT16_184 delay_INT16_184_2136 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2154:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x1_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:556:100
    .out   (_delay_INT16_184_2136_out)
  );
  delay_INT16_26 delay_INT16_26_2137 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2155:114
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:783:100
    .out   (_delay_INT16_26_2137_out)
  );
  delay_INT16_82 delay_INT16_82_2138 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2156:114
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x6_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1546:100
    .out   (_delay_INT16_82_2138_out)
  );
  delay_INT16_131 delay_INT16_131_2139 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2157:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_n_t6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:575:100
    .out   (_delay_INT16_131_2139_out)
  );
  delay_INT16_24 delay_INT16_24_2140 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2158:114
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x7_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:562:100
    .out   (_delay_INT16_24_2140_out)
  );
  delay_INT16_28 delay_INT16_28_2141 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2159:114
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x4_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:559:100
    .out   (_delay_INT16_28_2141_out)
  );
  delay_INT16_339 delay_INT16_339_2142 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2160:118
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x0_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:805:100
    .out   (_delay_INT16_339_2142_out)
  );
  delay_INT16_60 delay_INT16_60_2143 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2161:114
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x4_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:559:100
    .out   (_delay_INT16_60_2143_out)
  );
  delay_INT16_57 delay_INT16_57_2144 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2162:114
    .clock (clock),
    .reset (reset),
    .in    (_col_6_n_u7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1686:100
    .out   (_delay_INT16_57_2144_out)
  );
  delay_INT16_248 delay_INT16_248_2145 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2163:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_n_t3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:591:100
    .out   (_delay_INT16_248_2145_out)
  );
  delay_INT16_48 delay_INT16_48_2146 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2164:114
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x0_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:849:100
    .out   (_delay_INT16_48_2146_out)
  );
  delay_INT16_127 delay_INT16_127_2147 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2165:118
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:497:100
    .out   (_delay_INT16_127_2147_out)
  );
  delay_INT16_157 delay_INT16_157_2148 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2166:118
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:509:100
    .out   (_delay_INT16_157_2148_out)
  );
  delay_INT16_152 delay_INT16_152_2149 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2167:118
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:511:100
    .out   (_delay_INT16_152_2149_out)
  );
  delay_INT16_31 delay_INT16_31_2150 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2168:114
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x6_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:501:100
    .out   (_delay_INT16_31_2150_out)
  );
  delay_INT16_477 delay_INT16_477_2151 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2169:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x0_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1013:100
    .out   (_delay_INT16_477_2151_out)
  );
  delay_INT16_157 delay_INT16_157_2152 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2170:118
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x3_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:509:100
    .out   (_delay_INT16_157_2152_out)
  );
  delay_INT16_127 delay_INT16_127_2153 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2171:118
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x1_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:497:100
    .out   (_delay_INT16_127_2153_out)
  );
  delay_INT16_125 delay_INT16_125_2154 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2172:118
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:499:100
    .out   (_delay_INT16_125_2154_out)
  );
  delay_INT16_125 delay_INT16_125_2155 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2173:118
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x4_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:499:100
    .out   (_delay_INT16_125_2155_out)
  );
  delay_INT16_51 delay_INT16_51_2156 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2174:114
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1827:100
    .out   (_delay_INT16_51_2156_out)
  );
  delay_INT16_40 delay_INT16_40_2157 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2175:114
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:486:100
    .out   (_delay_INT16_40_2157_out)
  );
  delay_INT16_119 delay_INT16_119_2158 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2176:118
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1483:100
    .out   (_delay_INT16_119_2158_out)
  );
  delay_INT16_49 delay_INT16_49_2159 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2177:114
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:473:100
    .out   (_delay_INT16_49_2159_out)
  );
  delay_INT16_49 delay_INT16_49_2160 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2178:114
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x5_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:473:100
    .out   (_delay_INT16_49_2160_out)
  );
  delay_INT16_11 delay_INT16_11_2161 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2179:114
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:470:100
    .out   (_delay_INT16_11_2161_out)
  );
  delay_INT16_11 delay_INT16_11_2162 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2180:114
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x4_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:470:100
    .out   (_delay_INT16_11_2162_out)
  );
  delay_INT16_96 delay_INT16_96_2163 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2181:114
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x2_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:459:100
    .out   (_delay_INT16_96_2163_out)
  );
  delay_INT16_206 delay_INT16_206_2164 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2182:118
    .clock (clock),
    .reset (reset),
    .in    (_row_3_n_t7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:480:100
    .out   (_delay_INT16_206_2164_out)
  );
  delay_INT16_80 delay_INT16_80_2165 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2183:114
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x7_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1597:100
    .out   (_delay_INT16_80_2165_out)
  );
  delay_INT16_11 delay_INT16_11_2166 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2184:114
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x7_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:464:100
    .out   (_delay_INT16_11_2166_out)
  );
  delay_INT16_60 delay_INT16_60_2167 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2185:114
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x7_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:464:100
    .out   (_delay_INT16_60_2167_out)
  );
  delay_INT16_53 delay_INT16_53_2168 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2186:114
    .clock (clock),
    .reset (reset),
    .in    (_row_3_n_t5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:471:100
    .out   (_delay_INT16_53_2168_out)
  );
  delay_INT16_64 delay_INT16_64_2169 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2187:114
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x5_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:462:100
    .out   (_delay_INT16_64_2169_out)
  );
  delay_INT16_40 delay_INT16_40_2170 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2188:114
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x0_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:486:100
    .out   (_delay_INT16_40_2170_out)
  );
  delay_INT16_104 delay_INT16_104_2171 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2189:118
    .clock (clock),
    .reset (reset),
    .in    (_row_3_n_t4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:468:100
    .out   (_delay_INT16_104_2171_out)
  );
  delay_INT16_93 delay_INT16_93_2172 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2190:114
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x5_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:462:100
    .out   (_delay_INT16_93_2172_out)
  );
  delay_INT16_16 delay_INT16_16_2173 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2191:114
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1715:100
    .out   (_delay_INT16_16_2173_out)
  );
  delay_INT16_184 delay_INT16_184_2174 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2192:118
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x6_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:697:100
    .out   (_delay_INT16_184_2174_out)
  );
  delay_INT16_74 delay_INT16_74_2175 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2193:114
    .clock (clock),
    .reset (reset),
    .in    (_row_3_n_t6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:477:100
    .out   (_delay_INT16_74_2175_out)
  );
  delay_INT16_143 delay_INT16_143_2176 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2194:118
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:399:100
    .out   (_delay_INT16_143_2176_out)
  );
  delay_INT16_225 delay_INT16_225_2177 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2195:118
    .clock (clock),
    .reset (reset),
    .in    (_col_5_n_u3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1584:100
    .out   (_delay_INT16_225_2177_out)
  );
  delay_INT16_139 delay_INT16_139_2178 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2196:118
    .clock (clock),
    .reset (reset),
    .in    (_row_6_n_t6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:771:100
    .out   (_delay_INT16_139_2178_out)
  );
  delay_INT16_191 delay_INT16_191_2179 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2197:118
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:411:100
    .out   (_delay_INT16_191_2179_out)
  );
  delay_INT16_39 delay_INT16_39_2180 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2198:114
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:752:100
    .out   (_delay_INT16_39_2180_out)
  );
  delay_INT16_302 delay_INT16_302_2181 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2199:118
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:413:100
    .out   (_delay_INT16_302_2181_out)
  );
  delay_INT16_10 delay_INT16_10_2182 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2200:114
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x8_4_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:409:100
    .out   (_delay_INT16_10_2182_out)
  );
  delay_INT16_302 delay_INT16_302_2183 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2201:118
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x0_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:413:100
    .out   (_delay_INT16_302_2183_out)
  );
  delay_INT16_191 delay_INT16_191_2184 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2202:118
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x3_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:411:100
    .out   (_delay_INT16_191_2184_out)
  );
  delay_INT16_184 delay_INT16_184_2185 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2203:118
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:697:100
    .out   (_delay_INT16_184_2185_out)
  );
  delay_INT16_143 delay_INT16_143_2186 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2204:118
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x1_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:399:100
    .out   (_delay_INT16_143_2186_out)
  );
  delay_INT16_184 delay_INT16_184_2187 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2205:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:556:100
    .out   (_delay_INT16_184_2187_out)
  );
  delay_INT16_72 delay_INT16_72_2188 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2206:114
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:401:100
    .out   (_delay_INT16_72_2188_out)
  );
  delay_INT16_161 delay_INT16_161_2189 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2207:118
    .clock (clock),
    .reset (reset),
    .in    (_col_7_d_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1809:100
    .out   (_delay_INT16_161_2189_out)
  );
  delay_INT16_63 delay_INT16_63_2190 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2208:114
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:695:100
    .out   (_delay_INT16_63_2190_out)
  );
  delay_INT16_72 delay_INT16_72_2191 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2209:114
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x4_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:401:100
    .out   (_delay_INT16_72_2191_out)
  );
  delay_INT16_27 delay_INT16_27_2192 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2210:114
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:394:100
    .out   (_delay_INT16_27_2192_out)
  );
  delay_INT16_186 delay_INT16_186_2193 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2211:118
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x0_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1575:100
    .out   (_delay_INT16_186_2193_out)
  );
  delay_INT16_180 delay_INT16_180_2194 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2212:118
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x1_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:458:100
    .out   (_delay_INT16_180_2194_out)
  );
  delay_INT16_27 delay_INT16_27_2195 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2213:114
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x2_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:394:100
    .out   (_delay_INT16_27_2195_out)
  );
  delay_INT16_132 delay_INT16_132_2196 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2214:118
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x8_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:386:100
    .out   (_delay_INT16_132_2196_out)
  );
  delay_INT16_143 delay_INT16_143_2197 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2215:118
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:375:100
    .out   (_delay_INT16_143_2197_out)
  );
  delay_INT16_143 delay_INT16_143_2198 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2216:118
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x5_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:375:100
    .out   (_delay_INT16_143_2198_out)
  );
  delay_INT16_34 delay_INT16_34_2199 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2217:114
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:372:100
    .out   (_delay_INT16_34_2199_out)
  );
  delay_INT16_34 delay_INT16_34_2200 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2218:114
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x4_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:372:100
    .out   (_delay_INT16_34_2200_out)
  );
  delay_INT16_61 delay_INT16_61_2201 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2219:114
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x8_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1573:100
    .out   (_delay_INT16_61_2201_out)
  );
  delay_INT16_188 delay_INT16_188_2202 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2220:118
    .clock (clock),
    .reset (reset),
    .in    (_row_2_n_t3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:395:100
    .out   (_delay_INT16_188_2202_out)
  );
  delay_INT16_74 delay_INT16_74_2203 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2221:114
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x3_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:362:100
    .out   (_delay_INT16_74_2203_out)
  );
  delay_INT16_71 delay_INT16_71_2204 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2222:114
    .clock (clock),
    .reset (reset),
    .in    (_row_2_n_t2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:392:100
    .out   (_delay_INT16_71_2204_out)
  );
  delay_INT16_78 delay_INT16_78_2205 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2223:114
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x4_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1201:100
    .out   (_delay_INT16_78_2205_out)
  );
  delay_INT16_106 delay_INT16_106_2206 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2224:118
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x3_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:362:100
    .out   (_delay_INT16_106_2206_out)
  );
  delay_INT16_109 delay_INT16_109_2207 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2225:118
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:484:100
    .out   (_delay_INT16_109_2207_out)
  );
  delay_INT16_117 delay_INT16_117_2208 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2226:118
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:359:100
    .out   (_delay_INT16_117_2208_out)
  );
  delay_INT16_217 delay_INT16_217_2209 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2227:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_n_u4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:962:100
    .out   (_delay_INT16_217_2209_out)
  );
  delay_INT16_117 delay_INT16_117_2210 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2228:118
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x0_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:359:100
    .out   (_delay_INT16_117_2210_out)
  );
  delay_INT16_161 delay_INT16_161_2211 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2229:118
    .clock (clock),
    .reset (reset),
    .in    (_row_2_n_t7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:382:100
    .out   (_delay_INT16_161_2211_out)
  );
  delay_INT16_289 delay_INT16_289_2212 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2230:118
    .clock (clock),
    .reset (reset),
    .in    (_row_3_n_t2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:490:100
    .out   (_delay_INT16_289_2212_out)
  );
  delay_INT16_149 delay_INT16_149_2213 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2231:118
    .clock (clock),
    .reset (reset),
    .in    (_row_2_n_t6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:379:100
    .out   (_delay_INT16_149_2213_out)
  );
  delay_INT16_10 delay_INT16_10_2214 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2232:114
    .clock (clock),
    .reset (reset),
    .in    (_row_2_n_t4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:370:100
    .out   (_delay_INT16_10_2214_out)
  );
  delay_INT16_36 delay_INT16_36_2215 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2233:114
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x5_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:364:100
    .out   (_delay_INT16_36_2215_out)
  );
  delay_INT16_114 delay_INT16_114_2216 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2234:118
    .clock (clock),
    .reset (reset),
    .in    (_col_6_n_u6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1682:100
    .out   (_delay_INT16_114_2216_out)
  );
  delay_INT16_58 delay_INT16_58_2217 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2235:114
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x8_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:605:100
    .out   (_delay_INT16_58_2217_out)
  );
  delay_INT16_180 delay_INT16_180_2218 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2236:118
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:458:100
    .out   (_delay_INT16_180_2218_out)
  );
  delay_INT16_18 delay_INT16_18_2219 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2237:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:309:100
    .out   (_delay_INT16_18_2219_out)
  );
  delay_INT16_378 delay_INT16_378_2220 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2238:118
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x4_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1555:100
    .out   (_delay_INT16_378_2220_out)
  );
  delay_INT16_268 delay_INT16_268_2221 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2239:118
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:313:100
    .out   (_delay_INT16_268_2221_out)
  );
  delay_INT16_303 delay_INT16_303_2222 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2240:118
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:315:100
    .out   (_delay_INT16_303_2222_out)
  );
  delay_INT16_109 delay_INT16_109_2223 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2241:118
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x8_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:484:100
    .out   (_delay_INT16_109_2223_out)
  );
  delay_INT16_235 delay_INT16_235_2224 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2242:118
    .clock (clock),
    .reset (reset),
    .in    (_col_4_n_u5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1438:100
    .out   (_delay_INT16_235_2224_out)
  );
  delay_INT16_187 delay_INT16_187_2225 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2243:118
    .clock (clock),
    .reset (reset),
    .in    (_col_3_d_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1323:100
    .out   (_delay_INT16_187_2225_out)
  );
  delay_INT16_70 delay_INT16_70_2226 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2244:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x6_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:305:100
    .out   (_delay_INT16_70_2226_out)
  );
  delay_INT16_303 delay_INT16_303_2227 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2245:118
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x0_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:315:100
    .out   (_delay_INT16_303_2227_out)
  );
  delay_INT16_268 delay_INT16_268_2228 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2246:118
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x3_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:313:100
    .out   (_delay_INT16_268_2228_out)
  );
  delay_INT16_18 delay_INT16_18_2229 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2247:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x7_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:309:100
    .out   (_delay_INT16_18_2229_out)
  );
  delay_INT16_100 delay_INT16_100_2230 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2248:118
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x7_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1429:100
    .out   (_delay_INT16_100_2230_out)
  );
  delay_INT16_64 delay_INT16_64_2231 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2249:114
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x5_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1205:100
    .out   (_delay_INT16_64_2231_out)
  );
  delay_INT16_115 delay_INT16_115_2232 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2250:118
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:680:100
    .out   (_delay_INT16_115_2232_out)
  );
  delay_INT16_48 delay_INT16_48_2233 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2251:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:303:100
    .out   (_delay_INT16_48_2233_out)
  );
  delay_INT16_48 delay_INT16_48_2234 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2252:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x4_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:303:100
    .out   (_delay_INT16_48_2234_out)
  );
  delay_INT16_70 delay_INT16_70_2235 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2253:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:305:100
    .out   (_delay_INT16_70_2235_out)
  );
  delay_INT16_153 delay_INT16_153_2236 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2254:118
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:290:100
    .out   (_delay_INT16_153_2236_out)
  );
  delay_INT16_153 delay_INT16_153_2237 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2255:118
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x0_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:290:100
    .out   (_delay_INT16_153_2237_out)
  );
  delay_INT16_85 delay_INT16_85_2238 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2256:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:288:100
    .out   (_delay_INT16_85_2238_out)
  );
  delay_INT16_85 delay_INT16_85_2239 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2257:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x8_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:288:100
    .out   (_delay_INT16_85_2239_out)
  );
  delay_INT16_126 delay_INT16_126_2240 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2258:118
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:277:100
    .out   (_delay_INT16_126_2240_out)
  );
  delay_INT16_126 delay_INT16_126_2241 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2259:118
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x5_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:277:100
    .out   (_delay_INT16_126_2241_out)
  );
  delay_INT16_85 delay_INT16_85_2242 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2260:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:274:100
    .out   (_delay_INT16_85_2242_out)
  );
  delay_INT16_85 delay_INT16_85_2243 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2261:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x4_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:274:100
    .out   (_delay_INT16_85_2243_out)
  );
  delay_INT16_61 delay_INT16_61_2244 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2262:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_n_t3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:297:100
    .out   (_delay_INT16_61_2244_out)
  );
  delay_INT16_139 delay_INT16_139_2245 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2263:118
    .clock (clock),
    .reset (reset),
    .in    (_row_1_n_t2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:294:100
    .out   (_delay_INT16_139_2245_out)
  );
  delay_INT16_10 delay_INT16_10_2246 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2264:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x2_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:263:100
    .out   (_delay_INT16_10_2246_out)
  );
  delay_INT16_61 delay_INT16_61_2247 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2265:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:262:100
    .out   (_delay_INT16_61_2247_out)
  );
  delay_INT16_83 delay_INT16_83_2248 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2266:114
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1689:100
    .out   (_delay_INT16_83_2248_out)
  );
  delay_INT16_61 delay_INT16_61_2249 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2267:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x1_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:262:100
    .out   (_delay_INT16_61_2249_out)
  );
  delay_INT16_89 delay_INT16_89_2250 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2268:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_n_t7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:284:100
    .out   (_delay_INT16_89_2250_out)
  );
  delay_INT16_6 delay_INT16_6_2251 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2269:110
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x3_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:887:100
    .out   (_delay_INT16_6_2251_out)
  );
  delay_INT16_109 delay_INT16_109_2252 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2270:118
    .clock (clock),
    .reset (reset),
    .in    (_row_1_n_t6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:281:100
    .out   (_delay_INT16_109_2252_out)
  );
  delay_INT16_29 delay_INT16_29_2253 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2271:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x6_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:267:100
    .out   (_delay_INT16_29_2253_out)
  );
  delay_INT16_14 delay_INT16_14_2254 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2272:114
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1709:100
    .out   (_delay_INT16_14_2254_out)
  );
  delay_INT16_97 delay_INT16_97_2255 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2273:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_n_t5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:275:100
    .out   (_delay_INT16_97_2255_out)
  );
  delay_INT16_26 delay_INT16_26_2256 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2274:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_n_t4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:272:100
    .out   (_delay_INT16_26_2256_out)
  );
  delay_INT16_23 delay_INT16_23_2257 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2275:114
    .clock (clock),
    .reset (reset),
    .in    (_row_1_d_x5_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:266:100
    .out   (_delay_INT16_23_2257_out)
  );
  delay_INT16_80 delay_INT16_80_2258 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2276:114
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1597:100
    .out   (_delay_INT16_80_2258_out)
  );
  delay_INT16_72 delay_INT16_72_2259 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2277:114
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x3_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:558:100
    .out   (_delay_INT16_72_2259_out)
  );
  delay_INT16_20 delay_INT16_20_2260 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2278:114
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:203:100
    .out   (_delay_INT16_20_2260_out)
  );
  delay_INT16_206 delay_INT16_206_2261 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2279:118
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x3_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:215:100
    .out   (_delay_INT16_206_2261_out)
  );
  delay_INT16_162 delay_INT16_162_2262 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2280:118
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:217:100
    .out   (_delay_INT16_162_2262_out)
  );
  delay_INT16_49 delay_INT16_49_2263 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2281:114
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x6_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:207:100
    .out   (_delay_INT16_49_2263_out)
  );
  delay_INT16_162 delay_INT16_162_2264 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2282:118
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x0_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:217:100
    .out   (_delay_INT16_162_2264_out)
  );
  delay_INT16_225 delay_INT16_225_2265 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2283:118
    .clock (clock),
    .reset (reset),
    .in    (_col_7_n_u7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1804:100
    .out   (_delay_INT16_225_2265_out)
  );
  delay_INT16_206 delay_INT16_206_2266 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2284:118
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x3_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:215:100
    .out   (_delay_INT16_206_2266_out)
  );
  delay_INT16_20 delay_INT16_20_2267 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2285:114
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x1_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:203:100
    .out   (_delay_INT16_20_2267_out)
  );
  delay_INT16_75 delay_INT16_75_2268 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2286:114
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x3_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1233:100
    .out   (_delay_INT16_75_2268_out)
  );
  delay_INT16_89 delay_INT16_89_2269 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2287:114
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x4_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:205:100
    .out   (_delay_INT16_89_2269_out)
  );
  delay_INT16_89 delay_INT16_89_2270 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2288:114
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x4_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:205:100
    .out   (_delay_INT16_89_2270_out)
  );
  delay_INT16_106 delay_INT16_106_2271 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2289:118
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:192:100
    .out   (_delay_INT16_106_2271_out)
  );
  delay_INT16_120 delay_INT16_120_2272 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2290:118
    .clock (clock),
    .reset (reset),
    .in    (_row_6_d_x7_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:799:100
    .out   (_delay_INT16_120_2272_out)
  );
  delay_INT16_162 delay_INT16_162_2273 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2291:118
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:190:100
    .out   (_delay_INT16_162_2273_out)
  );
  delay_INT16_162 delay_INT16_162_2274 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2292:118
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x8_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:190:100
    .out   (_delay_INT16_162_2274_out)
  );
  delay_INT16_65 delay_INT16_65_2275 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2293:114
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:188:100
    .out   (_delay_INT16_65_2275_out)
  );
  delay_INT16_65 delay_INT16_65_2276 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2294:114
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x7_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:188:100
    .out   (_delay_INT16_65_2276_out)
  );
  delay_INT16_42 delay_INT16_42_2277 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2295:114
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:185:100
    .out   (_delay_INT16_42_2277_out)
  );
  delay_INT16_137 delay_INT16_137_2278 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2296:118
    .clock (clock),
    .reset (reset),
    .in    (_row_6_n_t4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:762:100
    .out   (_delay_INT16_137_2278_out)
  );
  delay_INT16_42 delay_INT16_42_2279 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2297:114
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x6_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:185:100
    .out   (_delay_INT16_42_2279_out)
  );
  delay_INT16_31 delay_INT16_31_2280 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2298:114
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:501:100
    .out   (_delay_INT16_31_2280_out)
  );
  delay_INT16_127 delay_INT16_127_2281 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2299:118
    .clock (clock),
    .reset (reset),
    .in    (_row_0_n_t3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:199:100
    .out   (_delay_INT16_127_2281_out)
  );
  delay_INT16_147 delay_INT16_147_2282 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2300:118
    .clock (clock),
    .reset (reset),
    .in    (_row_0_n_t2_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:196:100
    .out   (_delay_INT16_147_2282_out)
  );
  delay_INT16_27 delay_INT16_27_2283 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2301:114
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x2_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:165:100
    .out   (_delay_INT16_27_2283_out)
  );
  delay_INT16_350 delay_INT16_350_2284 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2302:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x0_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:609:100
    .out   (_delay_INT16_350_2284_out)
  );
  delay_INT16_100 delay_INT16_100_2285 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2303:118
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x2_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:165:100
    .out   (_delay_INT16_100_2285_out)
  );
  delay_INT16_245 delay_INT16_245_2286 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2304:118
    .clock (clock),
    .reset (reset),
    .in    (_col_7_n_u4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1788:100
    .out   (_delay_INT16_245_2286_out)
  );
  delay_INT16_29 delay_INT16_29_2287 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2305:114
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x1_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:164:100
    .out   (_delay_INT16_29_2287_out)
  );
  delay_INT16_93 delay_INT16_93_2288 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2306:114
    .clock (clock),
    .reset (reset),
    .in    (_row_0_n_t7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:186:100
    .out   (_delay_INT16_93_2288_out)
  );
  delay_INT16_15 delay_INT16_15_2289 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2307:114
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x7_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:170:100
    .out   (_delay_INT16_15_2289_out)
  );
  delay_INT16_171 delay_INT16_171_2290 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2308:118
    .clock (clock),
    .reset (reset),
    .in    (_row_0_n_t6_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:183:100
    .out   (_delay_INT16_171_2290_out)
  );
  delay_INT16_24 delay_INT16_24_2291 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2309:114
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x7_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:170:100
    .out   (_delay_INT16_24_2291_out)
  );
  delay_INT16_149 delay_INT16_149_2292 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2310:118
    .clock (clock),
    .reset (reset),
    .in    (_row_0_n_t5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:177:100
    .out   (_delay_INT16_149_2292_out)
  );
  delay_INT16_200 delay_INT16_200_2293 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2311:118
    .clock (clock),
    .reset (reset),
    .in    (_row_0_n_t4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:174:100
    .out   (_delay_INT16_200_2293_out)
  );
  delay_INT16_1 delay_INT16_1_2294 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2312:110
    .clock (clock),
    .reset (reset),
    .in    (_col_2_d_x6_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1192:100
    .out   (_delay_INT16_1_2294_out)
  );
  delay_INT16_45 delay_INT16_45_2295 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2313:114
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x4_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:167:100
    .out   (_delay_INT16_45_2295_out)
  );
  delay_INT16_7 delay_INT16_7_2296 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2314:110
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x6_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:365:100
    .out   (_delay_INT16_7_2296_out)
  );
  delay_INT16_106 delay_INT16_106_2297 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2315:118
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x0_1_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:192:100
    .out   (_delay_INT16_106_2297_out)
  );
  delay_INT16_108 delay_INT16_108_2298 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2316:118
    .clock (clock),
    .reset (reset),
    .in    (_row_3_n_t3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:493:100
    .out   (_delay_INT16_108_2298_out)
  );
  delay_INT16_268 delay_INT16_268_2299 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2317:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_n_t4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:566:100
    .out   (_delay_INT16_268_2299_out)
  );
  delay_INT16_61 delay_INT16_61_2300 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2318:114
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x8_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1573:100
    .out   (_delay_INT16_61_2300_out)
  );
  delay_INT16_29 delay_INT16_29_2301 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2319:114
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x1_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:164:100
    .out   (_delay_INT16_29_2301_out)
  );
  delay_INT16_2 delay_INT16_2_2302 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2320:110
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x1_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:881:100
    .out   (_delay_INT16_2_2302_out)
  );
  delay_INT16_104 delay_INT16_104_2303 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2321:118
    .clock (clock),
    .reset (reset),
    .in    (_row_2_n_t5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:373:100
    .out   (_delay_INT16_104_2303_out)
  );
  delay_INT16_193 delay_INT16_193_2304 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2322:118
    .clock (clock),
    .reset (reset),
    .in    (_col_3_n_u4_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1316:100
    .out   (_delay_INT16_193_2304_out)
  );
  delay_INT16_180 delay_INT16_180_2305 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2323:118
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x3_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1601:100
    .out   (_delay_INT16_180_2305_out)
  );
  delay_INT16_142 delay_INT16_142_2306 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2324:118
    .clock (clock),
    .reset (reset),
    .in    (_row_5_d_x1_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:693:100
    .out   (_delay_INT16_142_2306_out)
  );
  delay_INT16_152 delay_INT16_152_2307 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2325:118
    .clock (clock),
    .reset (reset),
    .in    (_row_3_d_x0_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:511:100
    .out   (_delay_INT16_152_2307_out)
  );
  delay_INT16_230 delay_INT16_230_2308 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2326:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_n_t5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:569:100
    .out   (_delay_INT16_230_2308_out)
  );
  delay_INT16_14 delay_INT16_14_2309 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2327:114
    .clock (clock),
    .reset (reset),
    .in    (_col_6_d_x4_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1709:100
    .out   (_delay_INT16_14_2309_out)
  );
  delay_INT16_306 delay_INT16_306_2310 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2328:118
    .clock (clock),
    .reset (reset),
    .in    (_col_7_n_u3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1820:100
    .out   (_delay_INT16_306_2310_out)
  );
  delay_INT16_158 delay_INT16_158_2311 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2329:118
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x3_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:953:100
    .out   (_delay_INT16_158_2311_out)
  );
  delay_INT16_10 delay_INT16_10_2312 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2330:114
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x8_4_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:409:100
    .out   (_delay_INT16_10_2312_out)
  );
  delay_INT16_119 delay_INT16_119_2313 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2331:118
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x3_2_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1483:100
    .out   (_delay_INT16_119_2313_out)
  );
  delay_INT16_378 delay_INT16_378_2314 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2332:118
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x5_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1559:100
    .out   (_delay_INT16_378_2314_out)
  );
  delay_INT16_34 delay_INT16_34_2315 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2333:114
    .clock (clock),
    .reset (reset),
    .in    (_col_0_d_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1003:100
    .out   (_delay_INT16_34_2315_out)
  );
  delay_INT16_19 delay_INT16_19_2316 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2334:114
    .clock (clock),
    .reset (reset),
    .in    (_row_7_d_x0_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:878:100
    .out   (_delay_INT16_19_2316_out)
  );
  delay_INT16_132 delay_INT16_132_2317 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2335:118
    .clock (clock),
    .reset (reset),
    .in    (_row_2_d_x8_3_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:386:100
    .out   (_delay_INT16_132_2317_out)
  );
  delay_INT16_234 delay_INT16_234_2318 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2336:118
    .clock (clock),
    .reset (reset),
    .in    (_row_4_n_t7_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:578:100
    .out   (_delay_INT16_234_2318_out)
  );
  delay_INT16_121 delay_INT16_121_2319 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2337:118
    .clock (clock),
    .reset (reset),
    .in    (_col_5_d_x0_0_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1540:100
    .out   (_delay_INT16_121_2319_out)
  );
  delay_INT16_23 delay_INT16_23_2320 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2338:114
    .clock (clock),
    .reset (reset),
    .in    (_col_6_n_u3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1702:100
    .out   (_delay_INT16_23_2320_out)
  );
  delay_INT16_6 delay_INT16_6_2321 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2339:110
    .clock (clock),
    .reset (reset),
    .in    (_col_4_d_x5_0_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1427:100
    .out   (_delay_INT16_6_2321_out)
  );
  delay_INT16_226 delay_INT16_226_2322 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2340:118
    .clock (clock),
    .reset (reset),
    .in    (_col_3_n_u3_1_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1348:100
    .out   (_delay_INT16_226_2322_out)
  );
  delay_INT16_49 delay_INT16_49_2323 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2341:114
    .clock (clock),
    .reset (reset),
    .in    (_row_0_d_x6_2_z),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:207:100
    .out   (_delay_INT16_49_2323_out)
  );
  delay_INT16_19 delay_INT16_19_2324 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2342:114
    .clock (clock),
    .reset (reset),
    .in    (_col_1_d_x4_3_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:1141:100
    .out   (_delay_INT16_19_2324_out)
  );
  delay_INT16_58 delay_INT16_58_2325 (	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:2343:114
    .clock (clock),
    .reset (reset),
    .in    (_row_4_d_x8_4_y),	// /home/nikita/Desktop/work/utopia/output/test/hil/idct/idctFir.mlir:605:100
    .out   (_delay_INT16_58_2325_out)
  );
endmodule

