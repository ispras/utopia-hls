// external module ADD_2x1

// external module MUL_2x1

// external module delay_fixed_16_0_1_11

// external module delay_fixed_16_0_1_22

// external module delay_fixed_16_0_1_25

// external module delay_fixed_16_0_1_34

// external module sink_1x0

// external module source_0x1

