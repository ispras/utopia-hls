module W2_add_W6(

    clock,
    reset,
    value);

output [15:0] value;
input clock;
input reset;
wire [15:0] value;
assign value = (2676+1108);
endmodule //W2_add_W6
