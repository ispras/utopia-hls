module IDCT(	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:11:5
  input         clock,
                reset,
  input  [15:0] source__dfc_wire_45__dfc_wire_45,
                source__dfc_wire_14__dfc_wire_45,
                source__dfc_wire_8__dfc_wire_45,
                source__dfc_wire_13__dfc_wire_45,
                source__dfc_wire_0__dfc_wire_45,
                source__dfc_wire_63__dfc_wire_45,
                source__dfc_wire_56__dfc_wire_45,
                source__dfc_wire_60__dfc_wire_45,
                source__dfc_wire_11__dfc_wire_45,
                source__dfc_wire_29__dfc_wire_45,
                source__dfc_wire_43__dfc_wire_45,
                source__dfc_wire_27__dfc_wire_45,
                source__dfc_wire_23__dfc_wire_45,
                source__dfc_wire_4__dfc_wire_45,
                source__dfc_wire_49__dfc_wire_45,
                source__dfc_wire_57__dfc_wire_45,
                source__dfc_wire_52__dfc_wire_45,
                source__dfc_wire_31__dfc_wire_45,
                source__dfc_wire_47__dfc_wire_45,
                source__dfc_wire_12__dfc_wire_45,
                source__dfc_wire_2__dfc_wire_45,
                source__dfc_wire_37__dfc_wire_45,
                source__dfc_wire_25__dfc_wire_45,
                source__dfc_wire_33__dfc_wire_45,
                source__dfc_wire_30__dfc_wire_45,
                source__dfc_wire_46__dfc_wire_45,
                source__dfc_wire_38__dfc_wire_45,
                source__dfc_wire_59__dfc_wire_45,
                source__dfc_wire_51__dfc_wire_45,
                source__dfc_wire_17__dfc_wire_45,
                source__dfc_wire_36__dfc_wire_45,
                source__dfc_wire_21__dfc_wire_45,
                source__dfc_wire_5__dfc_wire_45,
                source__dfc_wire_3__dfc_wire_45,
                source__dfc_wire_1__dfc_wire_45,
                source__dfc_wire_61__dfc_wire_45,
                source__dfc_wire_39__dfc_wire_45,
                source__dfc_wire_16__dfc_wire_45,
                source__dfc_wire_24__dfc_wire_45,
                source__dfc_wire_6__dfc_wire_45,
                source__dfc_wire_58__dfc_wire_45,
                source__dfc_wire_28__dfc_wire_45,
                source__dfc_wire_20__dfc_wire_45,
                source__dfc_wire_19__dfc_wire_45,
                source__dfc_wire_53__dfc_wire_45,
                source__dfc_wire_48__dfc_wire_45,
                source__dfc_wire_15__dfc_wire_45,
                source__dfc_wire_9__dfc_wire_45,
                source__dfc_wire_35__dfc_wire_45,
                source__dfc_wire_34__dfc_wire_45,
                source__dfc_wire_40__dfc_wire_45,
                source__dfc_wire_54__dfc_wire_45,
                source__dfc_wire_41__dfc_wire_45,
                source__dfc_wire_62__dfc_wire_45,
                source__dfc_wire_26__dfc_wire_45,
                source__dfc_wire_32__dfc_wire_45,
                source__dfc_wire_50__dfc_wire_45,
                source__dfc_wire_55__dfc_wire_45,
                source__dfc_wire_7__dfc_wire_45,
                source__dfc_wire_22__dfc_wire_45,
                source__dfc_wire_18__dfc_wire_45,
                source__dfc_wire_44__dfc_wire_45,
                source__dfc_wire_42__dfc_wire_45,
                source__dfc_wire_10__dfc_wire_45,
  output [15:0] sink__dfc_wire_4799__dfc_wire_4799,
                sink__dfc_wire_4777__dfc_wire_4799,
                sink__dfc_wire_4733__dfc_wire_4799,
                sink__dfc_wire_4711__dfc_wire_4799,
                sink__dfc_wire_4667__dfc_wire_4799,
                sink__dfc_wire_4369__dfc_wire_4799,
                sink__dfc_wire_4347__dfc_wire_4799,
                sink__dfc_wire_4303__dfc_wire_4799,
                sink__dfc_wire_4093__dfc_wire_4799,
                sink__dfc_wire_4049__dfc_wire_4799,
                sink__dfc_wire_4027__dfc_wire_4799,
                sink__dfc_wire_4005__dfc_wire_4799,
                sink__dfc_wire_3983__dfc_wire_4799,
                sink__dfc_wire_3961__dfc_wire_4799,
                sink__dfc_wire_3939__dfc_wire_4799,
                sink__dfc_wire_3707__dfc_wire_4799,
                sink__dfc_wire_3685__dfc_wire_4799,
                sink__dfc_wire_3597__dfc_wire_4799,
                sink__dfc_wire_3365__dfc_wire_4799,
                sink__dfc_wire_3321__dfc_wire_4799,
                sink__dfc_wire_3575__dfc_wire_4799,
                sink__dfc_wire_3277__dfc_wire_4799,
                sink__dfc_wire_3211__dfc_wire_4799,
                sink__dfc_wire_3343__dfc_wire_4799,
                sink__dfc_wire_2979__dfc_wire_4799,
                sink__dfc_wire_2913__dfc_wire_4799,
                sink__dfc_wire_3299__dfc_wire_4799,
                sink__dfc_wire_2637__dfc_wire_4799,
                sink__dfc_wire_2615__dfc_wire_4799,
                sink__dfc_wire_2593__dfc_wire_4799,
                sink__dfc_wire_2571__dfc_wire_4799,
                sink__dfc_wire_2549__dfc_wire_4799,
                sink__dfc_wire_2505__dfc_wire_4799,
                sink__dfc_wire_2483__dfc_wire_4799,
                sink__dfc_wire_3729__dfc_wire_4799,
                sink__dfc_wire_4689__dfc_wire_4799,
                sink__dfc_wire_2891__dfc_wire_4799,
                sink__dfc_wire_2163__dfc_wire_4799,
                sink__dfc_wire_3619__dfc_wire_4799,
                sink__dfc_wire_4755__dfc_wire_4799,
                sink__dfc_wire_4325__dfc_wire_4799,
                sink__dfc_wire_4071__dfc_wire_4799,
                sink__dfc_wire_4391__dfc_wire_4799,
                sink__dfc_wire_2251__dfc_wire_4799,
                sink__dfc_wire_2273__dfc_wire_4799,
                sink__dfc_wire_2957__dfc_wire_4799,
                sink__dfc_wire_3255__dfc_wire_4799,
                sink__dfc_wire_2185__dfc_wire_4799,
                sink__dfc_wire_2527__dfc_wire_4799,
                sink__dfc_wire_2935__dfc_wire_4799,
                sink__dfc_wire_4435__dfc_wire_4799,
                sink__dfc_wire_4457__dfc_wire_4799,
                sink__dfc_wire_2207__dfc_wire_4799,
                sink__dfc_wire_2869__dfc_wire_4799,
                sink__dfc_wire_2847__dfc_wire_4799,
                sink__dfc_wire_4413__dfc_wire_4799,
                sink__dfc_wire_2141__dfc_wire_4799,
                sink__dfc_wire_2229__dfc_wire_4799,
                sink__dfc_wire_2119__dfc_wire_4799,
                sink__dfc_wire_3233__dfc_wire_4799,
                sink__dfc_wire_3641__dfc_wire_4799,
                sink__dfc_wire_3001__dfc_wire_4799,
                sink__dfc_wire_4821__dfc_wire_4799,
                sink__dfc_wire_3663__dfc_wire_4799);

  wire [31:0] _delay_fixed_32_0_1_119_3245_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3263:146
  wire [31:0] _delay_fixed_32_0_1_12_3244_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3262:142
  wire [31:0] _delay_fixed_32_0_1_70_3243_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3261:142
  wire [31:0] _delay_fixed_32_0_1_34_3242_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3260:142
  wire [31:0] _delay_fixed_32_0_1_167_3241_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3259:146
  wire [31:0] _delay_fixed_32_0_1_1698_3240_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3258:150
  wire [31:0] _delay_fixed_32_0_1_55_3239_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3257:142
  wire [31:0] _delay_fixed_32_0_1_90_3238_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3256:142
  wire [31:0] _delay_fixed_32_0_1_1609_3237_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3255:150
  wire [31:0] _delay_fixed_32_0_1_93_3236_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3254:142
  wire [31:0] _delay_fixed_32_0_1_1715_3235_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3253:150
  wire        _delay_fixed_1_0_0_92_3234_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3252:138
  wire [31:0] _delay_fixed_32_0_1_140_3233_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3251:146
  wire [31:0] _delay_fixed_32_0_1_340_3232_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3250:146
  wire [31:0] _delay_fixed_32_0_1_230_3231_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3249:146
  wire [31:0] _delay_fixed_32_0_1_741_3230_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3248:146
  wire [31:0] _delay_fixed_32_0_1_246_3229_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3247:146
  wire [31:0] _delay_fixed_32_0_1_342_3228_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3246:146
  wire [31:0] _delay_fixed_32_0_1_72_3227_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3245:142
  wire [31:0] _delay_fixed_32_0_1_148_3226_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3244:146
  wire [31:0] _delay_fixed_32_0_1_23_3225_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3243:142
  wire [31:0] _delay_fixed_32_0_1_10_3224_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3242:142
  wire [31:0] _delay_fixed_32_0_1_280_3223_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3241:146
  wire [31:0] _delay_fixed_32_0_1_1411_3222_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3240:150
  wire [31:0] _delay_fixed_32_0_1_1417_3221_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3239:150
  wire [31:0] _delay_fixed_32_0_1_6_3220_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3238:138
  wire [31:0] _delay_fixed_32_0_1_5_3219_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3237:138
  wire [31:0] _delay_fixed_32_0_1_1377_3218_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3236:150
  wire [31:0] _delay_fixed_32_0_1_5_3217_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3235:138
  wire [31:0] _delay_fixed_32_0_1_1439_3216_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3234:150
  wire        _delay_fixed_1_0_0_15_3215_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3233:138
  wire [31:0] _delay_fixed_32_0_1_340_3214_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3232:146
  wire [31:0] _delay_fixed_32_0_1_1_3213_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3231:138
  wire [31:0] _delay_fixed_32_0_1_90_3212_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3230:142
  wire [31:0] _delay_fixed_32_0_1_130_3211_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3229:146
  wire [31:0] _delay_fixed_32_0_1_128_3210_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3228:146
  wire [31:0] _delay_fixed_32_0_1_188_3209_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3227:146
  wire [31:0] _delay_fixed_32_0_1_100_3208_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3226:146
  wire [31:0] _delay_fixed_32_0_1_85_3207_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3225:142
  wire [31:0] _delay_fixed_32_0_1_222_3206_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3224:146
  wire [31:0] _delay_fixed_32_0_1_157_3205_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3223:146
  wire [31:0] _delay_fixed_32_0_1_77_3204_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3222:142
  wire [31:0] _delay_fixed_32_0_1_905_3203_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3221:146
  wire [31:0] _delay_fixed_32_0_1_259_3202_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3220:146
  wire [31:0] _delay_fixed_32_0_1_11_3201_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3219:142
  wire [31:0] _delay_fixed_32_0_1_11_3200_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3218:142
  wire [31:0] _delay_fixed_32_0_1_1770_3199_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3217:150
  wire [31:0] _delay_fixed_32_0_1_1786_3198_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3216:150
  wire [31:0] _delay_fixed_32_0_1_16_3197_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3215:142
  wire [31:0] _delay_fixed_32_0_1_1736_3196_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3214:150
  wire [31:0] _delay_fixed_32_0_1_22_3195_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3213:142
  wire [31:0] _delay_fixed_32_0_1_1774_3194_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3212:150
  wire [31:0] _delay_fixed_32_0_1_19_3193_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3211:142
  wire [31:0] _delay_fixed_32_0_1_22_3192_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3210:142
  wire [31:0] _delay_fixed_32_0_1_178_3191_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3209:146
  wire [31:0] _delay_fixed_32_0_1_178_3190_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3208:146
  wire [31:0] _delay_fixed_32_0_1_205_3189_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3207:146
  wire [31:0] _delay_fixed_32_0_1_205_3188_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3206:146
  wire [31:0] _delay_fixed_32_0_1_1_3187_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3205:138
  wire [31:0] _delay_fixed_32_0_1_484_3186_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3204:146
  wire [31:0] _delay_fixed_32_0_1_566_3185_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3203:146
  wire [31:0] _delay_fixed_32_0_1_1_3184_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3202:138
  wire [31:0] _delay_fixed_32_0_1_461_3183_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3201:146
  wire [31:0] _delay_fixed_32_0_1_552_3182_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3200:146
  wire [31:0] _delay_fixed_32_0_1_46_3181_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3199:142
  wire [31:0] _delay_fixed_32_0_1_232_3180_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3198:146
  wire [31:0] _delay_fixed_32_0_1_139_3179_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3197:146
  wire [31:0] _delay_fixed_32_0_1_81_3178_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3196:142
  wire [31:0] _delay_fixed_32_0_1_81_3177_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3195:142
  wire [31:0] _delay_fixed_32_0_1_2274_3176_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3194:150
  wire        _delay_fixed_1_0_0_85_3175_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3193:138
  wire [31:0] _delay_fixed_32_0_1_139_3174_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3192:146
  wire [31:0] _delay_fixed_32_0_1_365_3173_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3191:146
  wire [31:0] _delay_fixed_32_0_1_232_3172_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3190:146
  wire [31:0] _delay_fixed_32_0_1_1987_3171_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3189:150
  wire [31:0] _delay_fixed_32_0_1_46_3170_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3188:142
  wire [31:0] _delay_fixed_32_0_1_1991_3169_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3187:150
  wire [31:0] _delay_fixed_32_0_1_4_3168_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3186:138
  wire [31:0] _delay_fixed_32_0_1_1953_3167_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3185:150
  wire [31:0] _delay_fixed_32_0_1_2006_3166_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3184:150
  wire        _delay_fixed_1_0_0_2_3165_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3183:134
  wire [31:0] _delay_fixed_32_0_1_156_3164_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3182:146
  wire [31:0] _delay_fixed_32_0_1_1796_3163_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3181:150
  wire [31:0] _delay_fixed_32_0_1_1835_3162_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3180:150
  wire [31:0] _delay_fixed_32_0_1_39_3161_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3179:142
  wire [31:0] _delay_fixed_32_0_1_1762_3160_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3178:150
  wire [31:0] _delay_fixed_32_0_1_1895_3159_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3177:150
  wire        _delay_fixed_1_0_0_52_3158_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3176:138
  wire [31:0] _delay_fixed_32_0_1_113_3157_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3175:146
  wire [31:0] _delay_fixed_32_0_1_156_3156_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3174:146
  wire [31:0] _delay_fixed_32_0_1_54_3155_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3173:142
  wire [31:0] _delay_fixed_32_0_1_73_3154_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3172:142
  wire [31:0] _delay_fixed_32_0_1_1713_3153_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3171:150
  wire [31:0] _delay_fixed_32_0_1_9_3152_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3170:138
  wire [31:0] _delay_fixed_32_0_1_1784_3151_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3169:150
  wire [31:0] _delay_fixed_32_0_1_71_3150_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3168:142
  wire [31:0] _delay_fixed_32_0_1_1679_3149_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3167:150
  wire [31:0] _delay_fixed_32_0_1_117_3148_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3166:146
  wire [31:0] _delay_fixed_32_0_1_1774_3147_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3165:150
  wire        _delay_fixed_1_0_0_30_3146_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3164:138
  wire [31:0] _delay_fixed_32_0_1_107_3145_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3163:146
  wire [31:0] _delay_fixed_32_0_1_27_3144_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3162:142
  wire [31:0] _delay_fixed_32_0_1_22_3143_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3161:142
  wire [31:0] _delay_fixed_32_0_1_178_3142_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3160:146
  wire [31:0] _delay_fixed_32_0_1_26_3141_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3159:142
  wire [31:0] _delay_fixed_32_0_1_98_3140_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3158:142
  wire [31:0] _delay_fixed_32_0_1_62_3139_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3157:142
  wire [31:0] _delay_fixed_32_0_1_138_3138_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3156:146
  wire [31:0] _delay_fixed_32_0_1_162_3137_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3155:146
  wire [31:0] _delay_fixed_32_0_1_162_3136_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3154:146
  wire [31:0] _delay_fixed_32_0_1_91_3135_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3153:142
  wire [31:0] _delay_fixed_32_0_1_190_3134_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3152:146
  wire [31:0] _delay_fixed_32_0_1_9_3133_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3151:138
  wire [31:0] _delay_fixed_32_0_1_172_3132_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3150:146
  wire [31:0] _delay_fixed_32_0_1_156_3131_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3149:146
  wire [31:0] _delay_fixed_32_0_1_98_3130_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3148:142
  wire [31:0] _delay_fixed_32_0_1_51_3129_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3147:142
  wire [31:0] _delay_fixed_32_0_1_51_3128_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3146:142
  wire [31:0] _delay_fixed_32_0_1_24_3127_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3145:142
  wire [31:0] _delay_fixed_32_0_1_24_3126_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3144:142
  wire [31:0] _delay_fixed_32_0_1_41_3125_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3143:142
  wire [31:0] _delay_fixed_32_0_1_41_3124_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3142:142
  wire [31:0] _delay_fixed_32_0_1_14_3123_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3141:142
  wire [31:0] _delay_fixed_32_0_1_14_3122_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3140:142
  wire [31:0] _delay_fixed_32_0_1_124_3121_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3139:146
  wire [31:0] _delay_fixed_32_0_1_486_3120_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3138:146
  wire [31:0] _delay_fixed_32_0_1_636_3119_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3137:146
  wire [31:0] _delay_fixed_32_0_1_124_3118_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3136:146
  wire [31:0] _delay_fixed_32_0_1_493_3117_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3135:146
  wire [31:0] _delay_fixed_32_0_1_624_3116_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3134:146
  wire [31:0] _delay_fixed_32_0_1_31_3115_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3133:142
  wire [31:0] _delay_fixed_32_0_1_461_3114_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3132:146
  wire [31:0] _delay_fixed_32_0_1_184_3113_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3131:146
  wire [31:0] _delay_fixed_32_0_1_110_3112_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3130:146
  wire [31:0] _delay_fixed_32_0_1_110_3111_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3129:146
  wire [31:0] _delay_fixed_32_0_1_184_3110_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3128:146
  wire [31:0] _delay_fixed_32_0_1_461_3109_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3127:146
  wire [31:0] _delay_fixed_32_0_1_31_3108_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3126:142
  wire [31:0] _delay_fixed_32_0_1_97_3107_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3125:142
  wire [31:0] _delay_fixed_32_0_1_122_3106_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3124:146
  wire [31:0] _delay_fixed_32_0_1_13_3105_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3123:142
  wire [31:0] _delay_fixed_32_0_1_143_3104_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3122:146
  wire [31:0] _delay_fixed_32_0_1_66_3103_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3121:142
  wire [31:0] _delay_fixed_32_0_1_225_3102_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3120:146
  wire [31:0] _delay_fixed_32_0_1_97_3101_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3119:142
  wire [31:0] _delay_fixed_32_0_1_212_3100_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3118:146
  wire [31:0] _delay_fixed_32_0_1_52_3099_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3117:142
  wire [31:0] _delay_fixed_32_0_1_256_3098_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3116:146
  wire [31:0] _delay_fixed_32_0_1_50_3097_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3115:142
  wire [31:0] _delay_fixed_32_0_1_146_3096_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3114:146
  wire [31:0] _delay_fixed_32_0_1_160_3095_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3113:146
  wire [31:0] _delay_fixed_32_0_1_270_3094_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3112:146
  wire [31:0] _delay_fixed_32_0_1_143_3093_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3111:146
  wire [31:0] _delay_fixed_32_0_1_53_3092_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3110:142
  wire [31:0] _delay_fixed_32_0_1_53_3091_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3109:142
  wire [31:0] _delay_fixed_32_0_1_216_3090_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3108:146
  wire [31:0] _delay_fixed_32_0_1_15_3089_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3107:142
  wire [31:0] _delay_fixed_32_0_1_83_3088_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3106:142
  wire [31:0] _delay_fixed_32_0_1_39_3087_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3105:142
  wire [31:0] _delay_fixed_32_0_1_17_3086_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3104:142
  wire [31:0] _delay_fixed_32_0_1_110_3085_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3103:146
  wire [31:0] _delay_fixed_32_0_1_110_3084_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3102:146
  wire [31:0] _delay_fixed_32_0_1_17_3083_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3101:142
  wire [31:0] _delay_fixed_32_0_1_33_3082_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3100:142
  wire [31:0] _delay_fixed_32_0_1_216_3081_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3099:146
  wire [31:0] _delay_fixed_32_0_1_37_3080_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3098:142
  wire [31:0] _delay_fixed_32_0_1_37_3079_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3097:142
  wire [31:0] _delay_fixed_32_0_1_365_3078_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3096:146
  wire [31:0] _delay_fixed_32_0_1_28_3077_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3095:142
  wire [31:0] _delay_fixed_32_0_1_28_3076_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3094:142
  wire [31:0] _delay_fixed_32_0_1_2076_3075_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3093:150
  wire [31:0] _delay_fixed_32_0_1_2139_3074_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3092:150
  wire [31:0] _delay_fixed_32_0_1_63_3073_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3091:142
  wire [31:0] _delay_fixed_32_0_1_47_3072_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3090:142
  wire [31:0] _delay_fixed_32_0_1_2042_3071_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3089:150
  wire [31:0] _delay_fixed_32_0_1_47_3070_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3088:142
  wire [31:0] _delay_fixed_32_0_1_2172_3069_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3087:150
  wire        _delay_fixed_1_0_0_60_3068_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3086:138
  wire [31:0] _delay_fixed_32_0_1_749_3067_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3085:146
  wire [31:0] _delay_fixed_32_0_1_1070_3066_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3084:150
  wire [31:0] _delay_fixed_32_0_1_1100_3065_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3083:150
  wire [31:0] _delay_fixed_32_0_1_51_3064_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3082:142
  wire [31:0] _delay_fixed_32_0_1_209_3063_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3081:146
  wire [31:0] _delay_fixed_32_0_1_1327_3062_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3080:150
  wire [31:0] _delay_fixed_32_0_1_51_3061_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3079:142
  wire [31:0] _delay_fixed_32_0_1_125_3060_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3078:146
  wire [31:0] _delay_fixed_32_0_1_1370_3059_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3077:150
  wire [31:0] _delay_fixed_32_0_1_43_3058_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3076:142
  wire [31:0] _delay_fixed_32_0_1_835_3057_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3075:146
  wire [31:0] _delay_fixed_32_0_1_1293_3056_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3074:150
  wire [31:0] _delay_fixed_32_0_1_218_3055_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3073:146
  wire [31:0] _delay_fixed_32_0_1_861_3054_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3072:146
  wire [31:0] _delay_fixed_32_0_1_1377_3053_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3071:150
  wire [31:0] _delay_fixed_32_0_1_26_3052_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3070:142
  wire [31:0] _delay_fixed_32_0_1_31_3051_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3069:142
  wire [31:0] _delay_fixed_32_0_1_386_3050_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3068:146
  wire [31:0] _delay_fixed_32_0_1_574_3049_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3067:146
  wire [31:0] _delay_fixed_32_0_1_346_3048_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3066:146
  wire [31:0] _delay_fixed_32_0_1_717_3047_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3065:146
  wire [31:0] _delay_fixed_32_0_1_126_3046_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3064:146
  wire [31:0] _delay_fixed_32_0_1_31_3045_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3063:142
  wire [31:0] _delay_fixed_32_0_1_126_3044_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3062:146
  wire [31:0] _delay_fixed_32_0_1_87_3043_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3061:142
  wire [31:0] _delay_fixed_32_0_1_1714_3042_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3060:150
  wire [31:0] _delay_fixed_32_0_1_634_3041_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3059:146
  wire [31:0] _delay_fixed_32_0_1_1099_3040_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3058:150
  wire [31:0] _delay_fixed_32_0_1_1783_3039_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3057:150
  wire [31:0] _delay_fixed_32_0_1_69_3038_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3056:142
  wire [31:0] _delay_fixed_32_0_1_778_3037_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3055:146
  wire [31:0] _delay_fixed_32_0_1_1076_3036_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3054:150
  wire [31:0] _delay_fixed_32_0_1_1680_3035_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3053:150
  wire [31:0] _delay_fixed_32_0_1_86_3034_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3052:142
  wire [31:0] _delay_fixed_32_0_1_983_3033_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3051:146
  wire [31:0] _delay_fixed_32_0_1_1825_3032_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3050:150
  wire        _delay_fixed_1_0_0_94_3031_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3049:138
  wire [31:0] _delay_fixed_32_0_1_822_3030_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3048:146
  wire [31:0] _delay_fixed_32_0_1_94_3029_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3047:142
  wire [31:0] _delay_fixed_32_0_1_787_3028_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3046:146
  wire [31:0] _delay_fixed_32_0_1_954_3027_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3045:146
  wire [31:0] _delay_fixed_32_0_1_136_3026_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3044:146
  wire [31:0] _delay_fixed_32_0_1_359_3025_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3043:146
  wire [31:0] _delay_fixed_32_0_1_1711_3024_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3042:150
  wire [31:0] _delay_fixed_32_0_1_1724_3023_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3041:150
  wire [31:0] _delay_fixed_32_0_1_13_3022_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3040:142
  wire [31:0] _delay_fixed_32_0_1_757_3021_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3039:146
  wire [31:0] _delay_fixed_32_0_1_1677_3020_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3038:150
  wire [31:0] _delay_fixed_32_0_1_399_3019_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3037:146
  wire [31:0] _delay_fixed_32_0_1_159_3018_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3036:146
  wire [31:0] _delay_fixed_32_0_1_1753_3017_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3035:150
  wire [31:0] _delay_fixed_32_0_1_9_3016_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3034:138
  wire [31:0] _delay_fixed_32_0_1_25_3015_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3033:142
  wire [31:0] _delay_fixed_32_0_1_25_3014_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3032:142
  wire [31:0] _delay_fixed_32_0_1_39_3013_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3031:142
  wire [31:0] _delay_fixed_32_0_1_225_3012_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3030:146
  wire [31:0] _delay_fixed_32_0_1_480_3011_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3029:146
  wire [31:0] _delay_fixed_32_0_1_225_3010_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3028:146
  wire [31:0] _delay_fixed_32_0_1_287_3009_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3027:146
  wire [31:0] _delay_fixed_32_0_1_1455_3008_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3026:150
  wire [31:0] _delay_fixed_32_0_1_1037_3007_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3025:150
  wire [31:0] _delay_fixed_32_0_1_1500_3006_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3024:150
  wire [31:0] _delay_fixed_32_0_1_45_3005_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3023:142
  wire [31:0] _delay_fixed_32_0_1_966_3004_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3022:146
  wire [31:0] _delay_fixed_32_0_1_1421_3003_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3021:150
  wire [31:0] _delay_fixed_32_0_1_206_3002_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3020:146
  wire [31:0] _delay_fixed_32_0_1_689_3001_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3019:146
  wire [31:0] _delay_fixed_32_0_1_1501_3000_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3018:150
  wire        _delay_fixed_1_0_0_25_2999_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3017:138
  wire [31:0] _delay_fixed_32_0_1_206_2998_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3016:146
  wire [31:0] _delay_fixed_32_0_1_90_2997_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3015:142
  wire [31:0] _delay_fixed_32_0_1_461_2996_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3014:146
  wire [31:0] _delay_fixed_32_0_1_130_2995_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3013:146
  wire [31:0] _delay_fixed_32_0_1_1032_2994_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3012:150
  wire [31:0] _delay_fixed_32_0_1_480_2993_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3011:146
  wire [31:0] _delay_fixed_32_0_1_99_2992_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3010:142
  wire [31:0] _delay_fixed_32_0_1_99_2991_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3009:142
  wire [31:0] _delay_fixed_32_0_1_4_2990_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3008:138
  wire [31:0] _delay_fixed_32_0_1_4_2989_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3007:138
  wire [31:0] _delay_fixed_32_0_1_399_2988_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3006:146
  wire [31:0] _delay_fixed_32_0_1_6_2987_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3005:138
  wire [31:0] _delay_fixed_32_0_1_1404_2986_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3004:150
  wire [31:0] _delay_fixed_32_0_1_70_2985_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3003:142
  wire [31:0] _delay_fixed_32_0_1_94_2984_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3002:142
  wire [31:0] _delay_fixed_32_0_1_1557_2983_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3001:150
  wire [31:0] _delay_fixed_32_0_1_70_2982_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3000:142
  wire [31:0] _delay_fixed_32_0_1_6_2981_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2999:138
  wire [31:0] _delay_fixed_32_0_1_1391_2980_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2998:150
  wire [31:0] _delay_fixed_32_0_1_1564_2979_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2997:150
  wire [31:0] _delay_fixed_32_0_1_190_2978_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2996:146
  wire [31:0] _delay_fixed_32_0_1_122_2977_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2995:146
  wire [31:0] _delay_fixed_32_0_1_54_2976_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2994:142
  wire [31:0] _delay_fixed_32_0_1_113_2975_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2993:146
  wire [31:0] _delay_fixed_32_0_1_44_2974_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2992:142
  wire [31:0] _delay_fixed_32_0_1_60_2973_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2991:142
  wire [31:0] _delay_fixed_32_0_1_142_2972_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2990:146
  wire [31:0] _delay_fixed_32_0_1_39_2971_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2989:142
  wire [31:0] _delay_fixed_32_0_1_76_2970_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2988:142
  wire [31:0] _delay_fixed_32_0_1_199_2969_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2987:146
  wire [31:0] _delay_fixed_32_0_1_43_2968_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2986:142
  wire [31:0] _delay_fixed_32_0_1_94_2967_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2985:142
  wire [31:0] _delay_fixed_32_0_1_25_2966_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2984:142
  wire [31:0] _delay_fixed_32_0_1_186_2965_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2983:146
  wire [31:0] _delay_fixed_32_0_1_12_2964_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2982:142
  wire [31:0] _delay_fixed_32_0_1_12_2963_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2981:142
  wire [31:0] _delay_fixed_32_0_1_72_2962_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2980:142
  wire [31:0] _delay_fixed_32_0_1_136_2961_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2979:146
  wire [31:0] _delay_fixed_32_0_1_44_2960_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2978:142
  wire [31:0] _delay_fixed_32_0_1_155_2959_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2977:146
  wire [31:0] _delay_fixed_32_0_1_28_2958_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2976:142
  wire [31:0] _delay_fixed_32_0_1_253_2957_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2975:146
  wire [31:0] _delay_fixed_32_0_1_15_2956_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2974:142
  wire [31:0] _delay_fixed_32_0_1_15_2955_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2973:142
  wire [31:0] _delay_fixed_32_0_1_16_2954_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2972:142
  wire [31:0] _delay_fixed_32_0_1_16_2953_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2971:142
  wire [31:0] _delay_fixed_32_0_1_14_2952_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2970:142
  wire [31:0] _delay_fixed_32_0_1_14_2951_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2969:142
  wire [31:0] _delay_fixed_32_0_1_87_2950_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2968:142
  wire [31:0] _delay_fixed_32_0_1_87_2949_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2967:142
  wire [31:0] _delay_fixed_32_0_1_46_2948_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2966:142
  wire [31:0] _delay_fixed_32_0_1_482_2947_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2965:146
  wire [31:0] _delay_fixed_32_0_1_625_2946_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2964:146
  wire [31:0] _delay_fixed_32_0_1_46_2945_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2963:142
  wire [31:0] _delay_fixed_32_0_1_456_2944_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2962:146
  wire [31:0] _delay_fixed_32_0_1_609_2943_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2961:146
  wire [31:0] _delay_fixed_32_0_1_55_2942_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2960:142
  wire [31:0] _delay_fixed_32_0_1_270_2941_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2959:146
  wire [31:0] _delay_fixed_32_0_1_55_2940_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2958:142
  wire [31:0] _delay_fixed_32_0_1_132_2939_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2957:146
  wire [31:0] _delay_fixed_32_0_1_10_2938_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2956:142
  wire [31:0] _delay_fixed_32_0_1_162_2937_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2955:146
  wire [31:0] _delay_fixed_32_0_1_75_2936_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2954:142
  wire [31:0] _delay_fixed_32_0_1_57_2935_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2953:142
  wire [31:0] _delay_fixed_32_0_1_166_2934_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2952:146
  wire [31:0] _delay_fixed_32_0_1_109_2933_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2951:146
  wire [31:0] _delay_fixed_32_0_1_30_2932_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2950:142
  wire [31:0] _delay_fixed_32_0_1_91_2931_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2949:142
  wire [31:0] _delay_fixed_32_0_1_7_2930_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2948:138
  wire [31:0] _delay_fixed_32_0_1_31_2929_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2947:142
  wire [31:0] _delay_fixed_32_0_1_21_2928_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2946:142
  wire [31:0] _delay_fixed_32_0_1_89_2927_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2945:142
  wire [31:0] _delay_fixed_32_0_1_11_2926_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2944:142
  wire [31:0] _delay_fixed_32_0_1_114_2925_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2943:146
  wire [31:0] _delay_fixed_32_0_1_10_2924_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2942:142
  wire [31:0] _delay_fixed_32_0_1_150_2923_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2941:146
  wire [31:0] _delay_fixed_32_0_1_79_2922_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2940:142
  wire [31:0] _delay_fixed_32_0_1_166_2921_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2939:146
  wire [31:0] _delay_fixed_32_0_1_4_2920_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2938:138
  wire [31:0] _delay_fixed_32_0_1_4_2919_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2937:138
  wire [31:0] _delay_fixed_32_0_1_66_2918_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2936:142
  wire [31:0] _delay_fixed_32_0_1_131_2917_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2935:146
  wire [31:0] _delay_fixed_32_0_1_81_2916_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2934:142
  wire [31:0] _delay_fixed_32_0_1_76_2915_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2933:142
  wire [31:0] _delay_fixed_32_0_1_71_2914_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2932:142
  wire [31:0] _delay_fixed_32_0_1_163_2913_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2931:146
  wire [31:0] _delay_fixed_32_0_1_72_2912_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2930:142
  wire [31:0] _delay_fixed_32_0_1_72_2911_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2929:142
  wire [31:0] _delay_fixed_32_0_1_40_2910_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2928:142
  wire [31:0] _delay_fixed_32_0_1_40_2909_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2927:142
  wire [31:0] _delay_fixed_32_0_1_45_2908_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2926:142
  wire [31:0] _delay_fixed_32_0_1_45_2907_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2925:142
  wire [31:0] _delay_fixed_32_0_1_47_2906_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2924:142
  wire [31:0] _delay_fixed_32_0_1_47_2905_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2923:142
  wire [31:0] _delay_fixed_32_0_1_103_2904_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2922:146
  wire [31:0] _delay_fixed_32_0_1_504_2903_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2921:146
  wire [31:0] _delay_fixed_32_0_1_605_2902_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2920:146
  wire [31:0] _delay_fixed_32_0_1_103_2901_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2919:146
  wire [31:0] _delay_fixed_32_0_1_473_2900_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2918:146
  wire [31:0] _delay_fixed_32_0_1_561_2899_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2917:146
  wire [31:0] _delay_fixed_32_0_1_57_2898_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2916:142
  wire [31:0] _delay_fixed_32_0_1_272_2897_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2915:146
  wire [31:0] _delay_fixed_32_0_1_212_2896_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2914:146
  wire [31:0] _delay_fixed_32_0_1_37_2895_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2913:142
  wire [31:0] _delay_fixed_32_0_1_37_2894_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2912:142
  wire [31:0] _delay_fixed_32_0_1_212_2893_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2911:146
  wire [31:0] _delay_fixed_32_0_1_272_2892_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2910:146
  wire [31:0] _delay_fixed_32_0_1_57_2891_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2909:142
  wire [31:0] _delay_fixed_32_0_1_131_2890_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2908:146
  wire [31:0] _delay_fixed_32_0_1_70_2889_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2907:142
  wire [31:0] _delay_fixed_32_0_1_145_2888_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2906:146
  wire [31:0] _delay_fixed_32_0_1_10_2887_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2905:142
  wire [31:0] _delay_fixed_32_0_1_103_2886_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2904:146
  wire [31:0] _delay_fixed_32_0_1_138_2885_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2903:146
  wire [31:0] _delay_fixed_32_0_1_3_2884_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2902:138
  wire [31:0] _delay_fixed_32_0_1_23_2883_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2901:142
  wire [31:0] _delay_fixed_32_0_1_23_2882_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2900:142
  wire [31:0] _delay_fixed_32_0_1_2_2881_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2899:138
  wire [31:0] _delay_fixed_32_0_1_177_2880_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2898:146
  wire [31:0] _delay_fixed_32_0_1_64_2879_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2897:142
  wire [31:0] _delay_fixed_32_0_1_110_2878_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2896:146
  wire [31:0] _delay_fixed_32_0_1_122_2877_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2895:146
  wire [31:0] _delay_fixed_32_0_1_95_2876_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2894:142
  wire [31:0] _delay_fixed_32_0_1_1_2875_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2893:138
  wire [31:0] _delay_fixed_32_0_1_1_2874_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2892:138
  wire [31:0] _delay_fixed_32_0_1_57_2873_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2891:142
  wire [31:0] _delay_fixed_32_0_1_57_2872_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2890:142
  wire [31:0] _delay_fixed_32_0_1_118_2871_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2889:146
  wire [31:0] _delay_fixed_32_0_1_118_2870_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2888:146
  wire [31:0] _delay_fixed_32_0_1_174_2869_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2887:146
  wire [31:0] _delay_fixed_32_0_1_174_2868_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2886:146
  wire [31:0] _delay_fixed_32_0_1_94_2867_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2885:142
  wire [31:0] _delay_fixed_32_0_1_497_2866_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2884:146
  wire [31:0] _delay_fixed_32_0_1_610_2865_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2883:146
  wire [31:0] _delay_fixed_32_0_1_94_2864_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2882:142
  wire [31:0] _delay_fixed_32_0_1_516_2863_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2881:146
  wire [31:0] _delay_fixed_32_0_1_670_2862_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2880:146
  wire [31:0] _delay_fixed_32_0_1_35_2861_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2879:142
  wire [31:0] _delay_fixed_32_0_1_134_2860_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2878:146
  wire [31:0] _delay_fixed_32_0_1_198_2859_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2877:146
  wire [31:0] _delay_fixed_32_0_1_73_2858_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2876:142
  wire [31:0] _delay_fixed_32_0_1_73_2857_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2875:142
  wire [31:0] _delay_fixed_32_0_1_198_2856_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2874:146
  wire [31:0] _delay_fixed_32_0_1_134_2855_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2873:146
  wire [31:0] _delay_fixed_32_0_1_35_2854_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2872:142
  wire [31:0] _delay_fixed_32_0_1_113_2853_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2871:146
  wire [31:0] _delay_fixed_32_0_1_73_2852_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2870:142
  wire [31:0] _delay_fixed_32_0_1_130_2851_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2869:146
  wire [31:0] _delay_fixed_32_0_1_202_2850_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2868:146
  wire [31:0] _delay_fixed_32_0_1_175_2849_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2867:146
  wire [31:0] _delay_fixed_32_0_1_24_2848_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2866:142
  wire [31:0] _delay_fixed_32_0_1_38_2847_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2865:142
  wire [31:0] _delay_fixed_32_0_1_146_2846_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2864:146
  wire [31:0] _delay_fixed_32_0_1_38_2845_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2863:142
  wire [31:0] _delay_fixed_32_0_1_30_2844_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2862:142
  wire [31:0] _delay_fixed_32_0_1_7_2843_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2861:138
  wire [31:0] _delay_fixed_32_0_1_29_2842_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2860:142
  wire [31:0] _delay_fixed_32_0_1_7_2841_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2859:138
  wire [31:0] _delay_fixed_32_0_1_164_2840_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2858:146
  wire [31:0] _delay_fixed_32_0_1_40_2839_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2857:142
  wire [31:0] _delay_fixed_32_0_1_70_2838_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2856:142
  wire [31:0] _delay_fixed_32_0_1_61_2837_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2855:142
  wire [31:0] _delay_fixed_32_0_1_70_2836_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2854:142
  wire [31:0] _delay_fixed_32_0_1_127_2835_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2853:146
  wire [31:0] _delay_fixed_32_0_1_11_2834_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2852:142
  wire [31:0] _delay_fixed_32_0_1_76_2833_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2851:142
  wire [31:0] _delay_fixed_32_0_1_76_2832_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2850:142
  wire [31:0] _delay_fixed_32_0_1_2_2831_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2849:138
  wire [31:0] _delay_fixed_32_0_1_2_2830_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2848:138
  wire [31:0] _delay_fixed_32_0_1_59_2829_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2847:142
  wire [31:0] _delay_fixed_32_0_1_1500_2828_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2846:150
  wire [31:0] _delay_fixed_32_0_1_129_2827_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2845:146
  wire [31:0] _delay_fixed_32_0_1_1646_2826_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2844:150
  wire [31:0] _delay_fixed_32_0_1_229_2825_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2843:146
  wire [31:0] _delay_fixed_32_0_1_1_2824_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2842:138
  wire [31:0] _delay_fixed_32_0_1_59_2823_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2841:142
  wire [31:0] _delay_fixed_32_0_1_1568_2822_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2840:150
  wire [31:0] _delay_fixed_32_0_1_247_2821_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2839:146
  wire [31:0] _delay_fixed_32_0_1_1685_2820_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2838:150
  wire [31:0] _delay_fixed_32_0_1_186_2819_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2837:146
  wire [31:0] _delay_fixed_32_0_1_132_2818_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2836:146
  wire [31:0] _delay_fixed_32_0_1_158_2817_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2835:146
  wire [31:0] _delay_fixed_32_0_1_30_2816_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2834:142
  wire [31:0] _delay_fixed_32_0_1_30_2815_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2833:142
  wire [31:0] _delay_fixed_32_0_1_1576_2814_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2832:150
  wire [31:0] _delay_fixed_32_0_1_1633_2813_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2831:150
  wire [31:0] _delay_fixed_32_0_1_57_2812_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2830:142
  wire [31:0] _delay_fixed_32_0_1_7_2811_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2829:138
  wire [31:0] _delay_fixed_32_0_1_1542_2810_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2828:150
  wire [31:0] _delay_fixed_32_0_1_7_2809_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2827:138
  wire [31:0] _delay_fixed_32_0_1_1657_2808_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2826:150
  wire        _delay_fixed_1_0_0_53_2807_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2825:138
  wire [31:0] _delay_fixed_32_0_1_258_2806_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2824:146
  wire [31:0] _delay_fixed_32_0_1_258_2805_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2823:146
  wire [31:0] _delay_fixed_32_0_1_440_2804_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2822:146
  wire [31:0] _delay_fixed_32_0_1_177_2803_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2821:146
  wire [31:0] _delay_fixed_32_0_1_1908_2802_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2820:150
  wire [31:0] _delay_fixed_32_0_1_177_2801_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2819:146
  wire [31:0] _delay_fixed_32_0_1_1959_2800_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2818:150
  wire [31:0] _delay_fixed_32_0_1_51_2799_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2817:142
  wire [31:0] _delay_fixed_32_0_1_1874_2798_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2816:150
  wire [31:0] _delay_fixed_32_0_1_1956_2797_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2815:150
  wire [31:0] _delay_fixed_32_0_1_19_2796_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2814:142
  wire [31:0] _delay_fixed_32_0_1_98_2795_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2813:142
  wire [31:0] _delay_fixed_32_0_1_417_2794_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2812:146
  wire [31:0] _delay_fixed_32_0_1_584_2793_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2811:146
  wire [31:0] _delay_fixed_32_0_1_445_2792_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2810:146
  wire [31:0] _delay_fixed_32_0_1_98_2791_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2809:142
  wire [31:0] _delay_fixed_32_0_1_442_2790_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2808:146
  wire [31:0] _delay_fixed_32_0_1_537_2789_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2807:146
  wire [31:0] _delay_fixed_32_0_1_1860_2788_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2806:150
  wire [31:0] _delay_fixed_32_0_1_1918_2787_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2805:150
  wire [31:0] _delay_fixed_32_0_1_58_2786_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2804:142
  wire [31:0] _delay_fixed_32_0_1_1826_2785_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2803:150
  wire [31:0] _delay_fixed_32_0_1_1912_2784_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2802:150
  wire        _delay_fixed_1_0_0_18_2783_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2801:138
  wire [31:0] _delay_fixed_32_0_1_90_2782_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2800:142
  wire [31:0] _delay_fixed_32_0_1_207_2781_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2799:146
  wire [31:0] _delay_fixed_32_0_1_65_2780_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2798:142
  wire [31:0] _delay_fixed_32_0_1_1693_2779_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2797:150
  wire [31:0] _delay_fixed_32_0_1_1758_2778_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2796:150
  wire [31:0] _delay_fixed_32_0_1_65_2777_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2795:142
  wire [31:0] _delay_fixed_32_0_1_1659_2776_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2794:150
  wire [31:0] _delay_fixed_32_0_1_1808_2775_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2793:150
  wire        _delay_fixed_1_0_0_79_2774_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2792:138
  wire [31:0] _delay_fixed_32_0_1_249_2773_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2791:146
  wire [31:0] _delay_fixed_32_0_1_207_2772_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2790:146
  wire [31:0] _delay_fixed_32_0_1_1727_2771_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2789:150
  wire [31:0] _delay_fixed_32_0_1_108_2770_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2788:146
  wire [31:0] _delay_fixed_32_0_1_1781_2769_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2787:150
  wire [31:0] _delay_fixed_32_0_1_54_2768_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2786:142
  wire [31:0] _delay_fixed_32_0_1_1693_2767_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2785:150
  wire [31:0] _delay_fixed_32_0_1_1806_2766_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2784:150
  wire        _delay_fixed_1_0_0_97_2765_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2783:138
  wire [31:0] _delay_fixed_32_0_1_108_2764_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2782:146
  wire [31:0] _delay_fixed_32_0_1_445_2763_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2781:146
  wire [31:0] _delay_fixed_32_0_1_249_2762_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2780:146
  wire [31:0] _delay_fixed_32_0_1_1936_2761_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2779:150
  wire [31:0] _delay_fixed_32_0_1_1968_2760_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2778:150
  wire [31:0] _delay_fixed_32_0_1_32_2759_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2777:142
  wire [31:0] _delay_fixed_32_0_1_65_2758_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2776:142
  wire [31:0] _delay_fixed_32_0_1_1902_2757_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2775:150
  wire [31:0] _delay_fixed_32_0_1_1980_2756_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2774:150
  wire        _delay_fixed_1_0_0_60_2755_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2773:138
  wire [31:0] _delay_fixed_32_0_1_90_2754_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2772:142
  wire [31:0] _delay_fixed_32_0_1_440_2753_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2771:146
  wire [31:0] _delay_fixed_32_0_1_1847_2752_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2770:150
  wire [31:0] _delay_fixed_32_0_1_1882_2751_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2769:150
  wire [31:0] _delay_fixed_32_0_1_35_2750_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2768:142
  wire [31:0] _delay_fixed_32_0_1_1813_2749_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2767:150
  wire [31:0] _delay_fixed_32_0_1_1899_2748_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2766:150
  wire        _delay_fixed_1_0_0_8_2747_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2765:134
  wire [31:0] _delay_fixed_32_0_1_158_2746_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2764:146
  wire [31:0] _delay_fixed_32_0_1_1583_2745_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2763:150
  wire [31:0] _delay_fixed_32_0_1_1624_2744_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2762:150
  wire [31:0] _delay_fixed_32_0_1_41_2743_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2761:142
  wire [31:0] _delay_fixed_32_0_1_134_2742_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2760:146
  wire [31:0] _delay_fixed_32_0_1_1549_2741_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2759:150
  wire [31:0] _delay_fixed_32_0_1_1597_2740_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2758:150
  wire        _delay_fixed_1_0_0_32_2739_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2757:138
  wire [31:0] _delay_fixed_32_0_1_13_2738_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2756:142
  wire [31:0] _delay_fixed_32_0_1_75_2737_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2755:142
  wire [31:0] _delay_fixed_32_0_1_4_2736_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2754:138
  wire [31:0] _delay_fixed_32_0_1_88_2735_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2753:142
  wire [31:0] _delay_fixed_32_0_1_53_2734_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2752:142
  wire [31:0] _delay_fixed_32_0_1_122_2733_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2751:146
  wire [31:0] _delay_fixed_32_0_1_82_2732_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2750:142
  wire [31:0] _delay_fixed_32_0_1_124_2731_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2749:146
  wire [31:0] _delay_fixed_32_0_1_765_2730_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2748:146
  wire [31:0] _delay_fixed_32_0_1_21_2729_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2747:142
  wire [31:0] _delay_fixed_32_0_1_131_2728_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2746:146
  wire [31:0] _delay_fixed_32_0_1_88_2727_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2745:142
  wire [31:0] _delay_fixed_32_0_1_119_2726_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2744:146
  wire [31:0] _delay_fixed_32_0_1_813_2725_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2743:146
  wire [31:0] _delay_fixed_32_0_1_17_2724_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2742:142
  wire [31:0] _delay_fixed_32_0_1_805_2723_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2741:146
  wire [31:0] _delay_fixed_32_0_1_647_2722_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2740:146
  wire [31:0] _delay_fixed_32_0_1_1560_2721_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2739:150
  wire [31:0] _delay_fixed_32_0_1_3_2720_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2738:138
  wire [31:0] _delay_fixed_32_0_1_1600_2719_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2737:150
  wire [31:0] _delay_fixed_32_0_1_40_2718_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2736:142
  wire [31:0] _delay_fixed_32_0_1_243_2717_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2735:146
  wire [31:0] _delay_fixed_32_0_1_3_2716_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2734:138
  wire [31:0] _delay_fixed_32_0_1_1526_2715_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2733:150
  wire [31:0] _delay_fixed_32_0_1_779_2714_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2732:146
  wire [31:0] _delay_fixed_32_0_1_1623_2713_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2731:150
  wire [31:0] _delay_fixed_32_0_1_53_2712_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2730:142
  wire [31:0] _delay_fixed_32_0_1_119_2711_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2729:146
  wire [31:0] _delay_fixed_32_0_1_80_2710_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2728:142
  wire [31:0] _delay_fixed_32_0_1_155_2709_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2727:146
  wire [31:0] _delay_fixed_32_0_1_98_2708_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2726:142
  wire [31:0] _delay_fixed_32_0_1_460_2707_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2725:146
  wire [31:0] _delay_fixed_32_0_1_131_2706_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2724:146
  wire [31:0] _delay_fixed_32_0_1_141_2705_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2723:146
  wire [31:0] _delay_fixed_32_0_1_808_2704_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2722:146
  wire [31:0] _delay_fixed_32_0_1_74_2703_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2721:142
  wire [31:0] _delay_fixed_32_0_1_742_2702_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2720:146
  wire [31:0] _delay_fixed_32_0_1_198_2701_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2719:146
  wire [31:0] _delay_fixed_32_0_1_1760_2700_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2718:150
  wire [31:0] _delay_fixed_32_0_1_725_2699_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2717:146
  wire [31:0] _delay_fixed_32_0_1_1787_2698_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2716:150
  wire [31:0] _delay_fixed_32_0_1_27_2697_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2715:142
  wire [31:0] _delay_fixed_32_0_1_1726_2696_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2714:150
  wire [31:0] _delay_fixed_32_0_1_176_2695_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2713:146
  wire [31:0] _delay_fixed_32_0_1_135_2694_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2712:146
  wire [31:0] _delay_fixed_32_0_1_1824_2693_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2711:150
  wire        _delay_fixed_1_0_0_36_2692_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2710:138
  wire [31:0] _delay_fixed_32_0_1_135_2691_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2709:146
  wire [31:0] _delay_fixed_32_0_1_652_2690_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2708:146
  wire [31:0] _delay_fixed_32_0_1_313_2689_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2707:146
  wire [31:0] _delay_fixed_32_0_1_1_2688_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2706:138
  wire [31:0] _delay_fixed_32_0_1_342_2687_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2705:146
  wire [31:0] _delay_fixed_32_0_1_1_2686_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2704:138
  wire [31:0] _delay_fixed_32_0_1_29_2685_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2703:142
  wire [31:0] _delay_fixed_32_0_1_1750_2684_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2702:150
  wire [31:0] _delay_fixed_32_0_1_29_2683_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2701:142
  wire [31:0] _delay_fixed_32_0_1_55_2682_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2700:142
  wire [31:0] _delay_fixed_32_0_1_1769_2681_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2699:150
  wire [31:0] _delay_fixed_32_0_1_19_2680_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2698:142
  wire [31:0] _delay_fixed_32_0_1_55_2679_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2697:142
  wire [31:0] _delay_fixed_32_0_1_1716_2678_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2696:150
  wire [31:0] _delay_fixed_32_0_1_1781_2677_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2695:150
  wire        _delay_fixed_1_0_0_27_2676_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2694:138
  wire [31:0] _delay_fixed_32_0_1_3_2675_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2693:138
  wire [31:0] _delay_fixed_32_0_1_769_2674_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2692:146
  wire [31:0] _delay_fixed_32_0_1_50_2673_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2691:142
  wire [31:0] _delay_fixed_32_0_1_658_2672_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2690:146
  wire [31:0] _delay_fixed_32_0_1_50_2671_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2689:142
  wire [31:0] _delay_fixed_32_0_1_673_2670_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2688:146
  wire [31:0] _delay_fixed_32_0_1_127_2669_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2687:146
  wire [31:0] _delay_fixed_32_0_1_195_2668_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2686:146
  wire [31:0] _delay_fixed_32_0_1_12_2667_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2685:142
  wire [31:0] _delay_fixed_32_0_1_472_2666_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2684:146
  wire [31:0] _delay_fixed_32_0_1_1433_2665_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2683:150
  wire [31:0] _delay_fixed_32_0_1_732_2664_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2682:146
  wire [31:0] _delay_fixed_32_0_1_552_2663_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2681:146
  wire [31:0] _delay_fixed_32_0_1_1529_2662_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2680:150
  wire [31:0] _delay_fixed_32_0_1_96_2661_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2679:142
  wire [31:0] _delay_fixed_32_0_1_174_2660_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2678:146
  wire [31:0] _delay_fixed_32_0_1_1399_2659_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2677:150
  wire [31:0] _delay_fixed_32_0_1_12_2658_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2676:142
  wire [31:0] _delay_fixed_32_0_1_1550_2657_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2675:150
  wire        _delay_fixed_1_0_0_108_2656_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2674:142
  wire [31:0] _delay_fixed_32_0_1_473_2655_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2673:146
  wire [31:0] _delay_fixed_32_0_1_622_2654_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2672:146
  wire [31:0] _delay_fixed_32_0_1_127_2653_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2671:146
  wire [31:0] _delay_fixed_32_0_1_3_2652_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2670:138
  wire [31:0] _delay_fixed_32_0_1_3_2651_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2669:138
  wire [31:0] _delay_fixed_32_0_1_1545_2650_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2668:150
  wire [31:0] _delay_fixed_32_0_1_85_2649_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2667:142
  wire [31:0] _delay_fixed_32_0_1_1571_2648_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2666:150
  wire [31:0] _delay_fixed_32_0_1_26_2647_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2665:142
  wire [31:0] _delay_fixed_32_0_1_75_2646_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2664:142
  wire [31:0] _delay_fixed_32_0_1_75_2645_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2663:142
  wire [31:0] _delay_fixed_32_0_1_235_2644_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2662:146
  wire [31:0] _delay_fixed_32_0_1_149_2643_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2661:146
  wire [31:0] _delay_fixed_32_0_1_235_2642_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2660:146
  wire [31:0] _delay_fixed_32_0_1_121_2641_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2659:146
  wire [31:0] _delay_fixed_32_0_1_121_2640_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2658:146
  wire [31:0] _delay_fixed_32_0_1_151_2639_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2657:146
  wire [31:0] _delay_fixed_32_0_1_24_2638_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2656:142
  wire [31:0] _delay_fixed_32_0_1_1238_2637_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2655:150
  wire [31:0] _delay_fixed_32_0_1_1362_2636_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2654:150
  wire [31:0] _delay_fixed_32_0_1_22_2635_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2653:142
  wire [31:0] _delay_fixed_32_0_1_24_2634_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2652:142
  wire [31:0] _delay_fixed_32_0_1_1277_2633_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2651:150
  wire [31:0] _delay_fixed_32_0_1_22_2632_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2650:142
  wire [31:0] _delay_fixed_32_0_1_1379_2631_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2649:150
  wire [31:0] _delay_fixed_32_0_1_1511_2630_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2648:150
  wire [31:0] _delay_fixed_32_0_1_1575_2629_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2647:150
  wire [31:0] _delay_fixed_32_0_1_11_2628_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2646:142
  wire [31:0] _delay_fixed_32_0_1_151_2627_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2645:146
  wire [31:0] _delay_fixed_32_0_1_342_2626_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2644:146
  wire [31:0] _delay_fixed_32_0_1_39_2625_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2643:142
  wire [31:0] _delay_fixed_32_0_1_149_2624_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2642:146
  wire [31:0] _delay_fixed_32_0_1_1736_2623_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2641:150
  wire [31:0] _delay_fixed_32_0_1_1488_2622_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2640:150
  wire [31:0] _delay_fixed_32_0_1_1758_2621_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2639:150
  wire [31:0] _delay_fixed_32_0_1_22_2620_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2638:142
  wire [31:0] _delay_fixed_32_0_1_1528_2619_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2637:150
  wire [31:0] _delay_fixed_32_0_1_40_2618_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2636:142
  wire [31:0] _delay_fixed_32_0_1_85_2617_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2635:142
  wire [31:0] _delay_fixed_32_0_1_1702_2616_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2634:150
  wire [31:0] _delay_fixed_32_0_1_1454_2615_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2633:150
  wire [31:0] _delay_fixed_32_0_1_1758_2614_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2632:150
  wire [31:0] _delay_fixed_32_0_1_33_2613_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2631:142
  wire [31:0] _delay_fixed_32_0_1_1575_2612_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2630:150
  wire        _delay_fixed_1_0_0_52_2611_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2629:138
  wire [31:0] _delay_fixed_32_0_1_460_2610_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2628:146
  wire [31:0] _delay_fixed_32_0_1_342_2609_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2627:146
  wire [31:0] _delay_fixed_32_0_1_1915_2608_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2626:150
  wire [31:0] _delay_fixed_32_0_1_1956_2607_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2625:150
  wire [31:0] _delay_fixed_32_0_1_41_2606_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2624:142
  wire [31:0] _delay_fixed_32_0_1_1881_2605_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2623:150
  wire [31:0] _delay_fixed_32_0_1_1643_2604_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2622:150
  wire [31:0] _delay_fixed_32_0_1_1963_2603_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2621:150
  wire        _delay_fixed_1_0_0_53_2602_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2620:138
  wire [31:0] _delay_fixed_32_0_1_1672_2601_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2619:150
  wire [31:0] _delay_fixed_32_0_1_29_2600_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2618:142
  wire [31:0] _delay_fixed_32_0_1_1609_2599_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2617:150
  wire [31:0] _delay_fixed_32_0_1_190_2598_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2616:146
  wire [31:0] _delay_fixed_32_0_1_1702_2597_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2615:150
  wire [31:0] _delay_fixed_32_0_1_62_2596_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2614:142
  wire [31:0] _delay_fixed_32_0_1_825_2595_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2613:146
  wire [31:0] _delay_fixed_32_0_1_1604_2594_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2612:150
  wire [31:0] _delay_fixed_32_0_1_1651_2593_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2611:150
  wire [31:0] _delay_fixed_32_0_1_47_2592_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2610:142
  wire [31:0] _delay_fixed_32_0_1_346_2591_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2609:146
  wire [31:0] _delay_fixed_32_0_1_1570_2590_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2608:150
  wire [31:0] _delay_fixed_32_0_1_41_2589_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2607:142
  wire [31:0] _delay_fixed_32_0_1_1666_2588_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2606:150
  wire [31:0] _delay_fixed_32_0_1_13_2587_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2605:142
  wire [31:0] _delay_fixed_32_0_1_744_2586_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2604:146
  wire [31:0] _delay_fixed_32_0_1_1692_2585_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2603:150
  wire [31:0] _delay_fixed_32_0_1_1658_2584_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2602:150
  wire [31:0] _delay_fixed_32_0_1_706_2583_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2601:146
  wire [31:0] _delay_fixed_32_0_1_1741_2582_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2600:150
  wire [31:0] _delay_fixed_32_0_1_19_2581_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2599:142
  wire [31:0] _delay_fixed_32_0_1_689_2580_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2598:146
  wire [31:0] _delay_fixed_32_0_1_60_2579_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2597:142
  wire [31:0] _delay_fixed_32_0_1_24_2578_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2596:142
  wire [31:0] _delay_fixed_32_0_1_692_2577_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2595:146
  wire [31:0] _delay_fixed_32_0_1_125_2576_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2594:146
  wire [31:0] _delay_fixed_32_0_1_1419_2575_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2593:150
  wire [31:0] _delay_fixed_32_0_1_1021_2574_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2592:150
  wire [31:0] _delay_fixed_32_0_1_1434_2573_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2591:150
  wire [31:0] _delay_fixed_32_0_1_15_2572_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2590:142
  wire [31:0] _delay_fixed_32_0_1_1385_2571_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2589:150
  wire [31:0] _delay_fixed_32_0_1_28_2570_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2588:142
  wire [31:0] _delay_fixed_32_0_1_1424_2569_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2587:150
  wire [31:0] _delay_fixed_32_0_1_6_2568_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2586:138
  wire [31:0] _delay_fixed_32_0_1_913_2567_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2585:146
  wire [31:0] _delay_fixed_32_0_1_283_2566_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2584:146
  wire [31:0] _delay_fixed_32_0_1_842_2565_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2583:146
  wire [31:0] _delay_fixed_32_0_1_1147_2564_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2582:150
  wire [31:0] _delay_fixed_32_0_1_24_2563_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2581:142
  wire [31:0] _delay_fixed_32_0_1_1715_2562_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2580:150
  wire [31:0] _delay_fixed_32_0_1_23_2561_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2579:142
  wire [31:0] _delay_fixed_32_0_1_256_2560_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2578:146
  wire [31:0] _delay_fixed_32_0_1_256_2559_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2577:146
  wire [31:0] _delay_fixed_32_0_1_226_2558_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2576:146
  wire [31:0] _delay_fixed_32_0_1_226_2557_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2575:146
  wire [31:0] _delay_fixed_32_0_1_80_2556_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2574:142
  wire [31:0] _delay_fixed_32_0_1_1728_2555_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2573:150
  wire [31:0] _delay_fixed_32_0_1_1838_2554_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2572:150
  wire [31:0] _delay_fixed_32_0_1_80_2553_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2571:142
  wire [31:0] _delay_fixed_32_0_1_1732_2552_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2570:150
  wire [31:0] _delay_fixed_32_0_1_1811_2551_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2569:150
  wire [31:0] _delay_fixed_32_0_1_59_2550_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2568:142
  wire [31:0] _delay_fixed_32_0_1_1747_2549_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2567:150
  wire [31:0] _delay_fixed_32_0_1_1786_2548_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2566:150
  wire [31:0] _delay_fixed_32_0_1_39_2547_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2565:142
  wire [31:0] _delay_fixed_32_0_1_1713_2546_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2564:150
  wire [31:0] _delay_fixed_32_0_1_1807_2545_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2563:150
  wire        _delay_fixed_1_0_0_75_2544_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2562:138
  wire [31:0] _delay_fixed_32_0_1_478_2543_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2561:146
  wire [31:0] _delay_fixed_32_0_1_2173_2542_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2560:150
  wire [31:0] _delay_fixed_32_0_1_2262_2541_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2559:150
  wire [31:0] _delay_fixed_32_0_1_89_2540_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2558:142
  wire [31:0] _delay_fixed_32_0_1_2139_2539_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2557:150
  wire [31:0] _delay_fixed_32_0_1_478_2538_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2556:146
  wire [31:0] _delay_fixed_32_0_1_2078_2537_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2555:150
  wire [31:0] _delay_fixed_32_0_1_2085_2536_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2554:150
  wire [31:0] _delay_fixed_32_0_1_7_2535_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2553:138
  wire [31:0] _delay_fixed_32_0_1_2044_2534_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2552:150
  wire [31:0] _delay_fixed_32_0_1_2086_2533_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2551:150
  wire        _delay_fixed_1_0_0_9_2532_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2550:134
  wire [31:0] _delay_fixed_32_0_1_59_2531_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2549:142
  wire [31:0] _delay_fixed_32_0_1_1678_2530_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2548:150
  wire [31:0] _delay_fixed_32_0_1_1717_2529_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2547:150
  wire [31:0] _delay_fixed_32_0_1_39_2528_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2546:142
  wire [31:0] _delay_fixed_32_0_1_1644_2527_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2545:150
  wire [31:0] _delay_fixed_32_0_1_1777_2526_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2544:150
  wire        _delay_fixed_1_0_0_95_2525_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2543:138
  wire [31:0] _delay_fixed_32_0_1_915_2524_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2542:146
  wire [31:0] _delay_fixed_32_0_1_155_2523_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2541:146
  wire [31:0] _delay_fixed_32_0_1_1014_2522_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2540:150
  wire [31:0] _delay_fixed_32_0_1_983_2521_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2539:146
  wire [31:0] _delay_fixed_32_0_1_781_2520_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2538:146
  wire [31:0] _delay_fixed_32_0_1_295_2519_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2537:146
  wire [31:0] _delay_fixed_32_0_1_980_2518_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2536:146
  wire [31:0] _delay_fixed_32_0_1_138_2517_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2535:146
  wire [31:0] _delay_fixed_32_0_1_73_2516_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2534:142
  wire [31:0] _delay_fixed_32_0_1_1032_2515_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2533:150
  wire [31:0] _delay_fixed_32_0_1_1009_2514_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2532:150
  wire [31:0] _delay_fixed_32_0_1_920_2513_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2531:146
  wire [31:0] _delay_fixed_32_0_1_122_2512_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2530:146
  wire [31:0] _delay_fixed_32_0_1_7_2511_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2529:138
  wire [31:0] _delay_fixed_32_0_1_1062_2510_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2528:150
  wire [31:0] _delay_fixed_32_0_1_986_2509_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2527:146
  wire [31:0] _delay_fixed_32_0_1_994_2508_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2526:146
  wire [31:0] _delay_fixed_32_0_1_123_2507_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2525:146
  wire [31:0] _delay_fixed_32_0_1_1043_2506_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2524:150
  wire [31:0] _delay_fixed_32_0_1_167_2505_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2523:146
  wire [31:0] _delay_fixed_32_0_1_1_2504_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2522:138
  wire [31:0] _delay_fixed_32_0_1_1_2503_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2521:138
  wire [31:0] _delay_fixed_32_0_1_25_2502_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2520:142
  wire [31:0] _delay_fixed_32_0_1_25_2501_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2519:142
  wire [31:0] _delay_fixed_32_0_1_270_2500_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2518:146
  wire [31:0] _delay_fixed_32_0_1_270_2499_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2517:146
  wire [31:0] _delay_fixed_32_0_1_172_2498_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2516:146
  wire [31:0] _delay_fixed_32_0_1_172_2497_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2515:146
  wire [31:0] _delay_fixed_32_0_1_111_2496_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2514:146
  wire [31:0] _delay_fixed_32_0_1_1578_2495_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2513:150
  wire [31:0] _delay_fixed_32_0_1_1687_2494_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2512:150
  wire [31:0] _delay_fixed_32_0_1_111_2493_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2511:146
  wire [31:0] _delay_fixed_32_0_1_1556_2492_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2510:150
  wire [31:0] _delay_fixed_32_0_1_1679_2491_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2509:150
  wire [31:0] _delay_fixed_32_0_1_102_2490_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2508:146
  wire [31:0] _delay_fixed_32_0_1_1726_2489_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2507:150
  wire [31:0] _delay_fixed_32_0_1_1818_2488_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2506:150
  wire [31:0] _delay_fixed_32_0_1_92_2487_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2505:142
  wire [31:0] _delay_fixed_32_0_1_1692_2486_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2504:150
  wire [31:0] _delay_fixed_32_0_1_1798_2485_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2503:150
  wire        _delay_fixed_1_0_0_13_2484_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2502:138
  wire [31:0] _delay_fixed_32_0_1_295_2483_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2501:146
  wire [31:0] _delay_fixed_32_0_1_1826_2482_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2500:150
  wire [31:0] _delay_fixed_32_0_1_1827_2481_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2499:150
  wire [31:0] _delay_fixed_32_0_1_1_2480_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2498:138
  wire [31:0] _delay_fixed_32_0_1_1792_2479_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2497:150
  wire [31:0] _delay_fixed_32_0_1_1876_2478_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2496:150
  wire        _delay_fixed_1_0_0_81_2477_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2495:138
  wire [31:0] _delay_fixed_32_0_1_356_2476_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2494:146
  wire [31:0] _delay_fixed_32_0_1_1825_2475_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2493:150
  wire [31:0] _delay_fixed_32_0_1_1869_2474_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2492:150
  wire [31:0] _delay_fixed_32_0_1_44_2473_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2491:142
  wire [31:0] _delay_fixed_32_0_1_1791_2472_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2490:150
  wire [31:0] _delay_fixed_32_0_1_1918_2471_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2489:150
  wire        _delay_fixed_1_0_0_80_2470_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2488:138
  wire [31:0] _delay_fixed_32_0_1_103_2469_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2487:146
  wire [31:0] _delay_fixed_32_0_1_1636_2468_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2486:150
  wire [31:0] _delay_fixed_32_0_1_1721_2467_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2485:150
  wire [31:0] _delay_fixed_32_0_1_85_2466_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2484:142
  wire [31:0] _delay_fixed_32_0_1_1602_2465_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2483:150
  wire [31:0] _delay_fixed_32_0_1_1759_2464_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2482:150
  wire        _delay_fixed_1_0_0_76_2463_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2481:138
  wire [31:0] _delay_fixed_32_0_1_103_2462_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2480:146
  wire [31:0] _delay_fixed_32_0_1_1722_2461_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2479:150
  wire [31:0] _delay_fixed_32_0_1_1761_2460_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2478:150
  wire [31:0] _delay_fixed_32_0_1_39_2459_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2477:142
  wire [31:0] _delay_fixed_32_0_1_1688_2458_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2476:150
  wire [31:0] _delay_fixed_32_0_1_1774_2457_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2475:150
  wire        _delay_fixed_1_0_0_7_2456_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2474:134
  wire [31:0] _delay_fixed_32_0_1_356_2455_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2473:146
  wire [31:0] _delay_fixed_32_0_1_1880_2454_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2472:150
  wire [31:0] _delay_fixed_32_0_1_1930_2453_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2471:150
  wire [31:0] _delay_fixed_32_0_1_50_2452_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2470:142
  wire [31:0] _delay_fixed_32_0_1_1846_2451_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2469:150
  wire [31:0] _delay_fixed_32_0_1_1941_2450_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2468:150
  wire        _delay_fixed_1_0_0_20_2449_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2467:138
  wire [31:0] _delay_fixed_32_0_1_295_2448_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2466:146
  wire [31:0] _delay_fixed_32_0_1_1915_2447_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2465:150
  wire [31:0] _delay_fixed_32_0_1_1972_2446_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2464:150
  wire [31:0] _delay_fixed_32_0_1_57_2445_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2463:142
  wire [31:0] _delay_fixed_32_0_1_1881_2444_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2462:150
  wire [31:0] _delay_fixed_32_0_1_2017_2443_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2461:150
  wire        _delay_fixed_1_0_0_75_2442_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2460:138
  wire [31:0] _delay_fixed_32_0_1_102_2441_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2459:146
  wire [31:0] _delay_fixed_32_0_1_1761_2440_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2458:150
  wire [31:0] _delay_fixed_32_0_1_1788_2439_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2457:150
  wire [31:0] _delay_fixed_32_0_1_27_2438_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2456:142
  wire [31:0] _delay_fixed_32_0_1_1727_2437_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2455:150
  wire [31:0] _delay_fixed_32_0_1_1775_2436_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2454:150
  wire        _delay_fixed_1_0_0_13_2435_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2453:138
  wire [31:0] _delay_fixed_32_0_1_835_2434_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2452:146
  wire [31:0] _delay_fixed_32_0_1_3_2433_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2451:138
  wire [31:0] _delay_fixed_32_0_1_744_2432_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2450:146
  wire [31:0] _delay_fixed_32_0_1_711_2431_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2449:146
  wire [31:0] _delay_fixed_32_0_1_729_2430_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2448:146
  wire [31:0] _delay_fixed_32_0_1_80_2429_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2447:142
  wire [31:0] _delay_fixed_32_0_1_776_2428_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2446:146
  wire [31:0] _delay_fixed_32_0_1_36_2427_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2445:142
  wire [31:0] _delay_fixed_32_0_1_9_2426_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2444:138
  wire [31:0] _delay_fixed_32_0_1_781_2425_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2443:146
  wire [31:0] _delay_fixed_32_0_1_678_2424_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2442:146
  wire [31:0] _delay_fixed_32_0_1_670_2423_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2441:146
  wire [31:0] _delay_fixed_32_0_1_130_2422_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2440:146
  wire [31:0] _delay_fixed_32_0_1_719_2421_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2439:146
  wire [31:0] _delay_fixed_32_0_1_71_2420_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2438:142
  wire [31:0] _delay_fixed_32_0_1_12_2419_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2437:142
  wire [31:0] _delay_fixed_32_0_1_12_2418_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2436:142
  wire [31:0] _delay_fixed_32_0_1_161_2417_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2435:146
  wire [31:0] _delay_fixed_32_0_1_869_2416_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2434:146
  wire [31:0] _delay_fixed_32_0_1_768_2415_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2433:146
  wire [31:0] _delay_fixed_32_0_1_622_2414_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2432:146
  wire [31:0] _delay_fixed_32_0_1_341_2413_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2431:146
  wire [31:0] _delay_fixed_32_0_1_839_2412_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2430:146
  wire [31:0] _delay_fixed_32_0_1_175_2411_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2429:146
  wire [31:0] _delay_fixed_32_0_1_11_2410_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2428:142
  wire [31:0] _delay_fixed_32_0_1_11_2409_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2427:142
  wire [31:0] _delay_fixed_32_0_1_39_2408_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2426:142
  wire [31:0] _delay_fixed_32_0_1_39_2407_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2425:142
  wire [31:0] _delay_fixed_32_0_1_169_2406_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2424:146
  wire [31:0] _delay_fixed_32_0_1_169_2405_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2423:146
  wire [31:0] _delay_fixed_32_0_1_288_2404_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2422:146
  wire [31:0] _delay_fixed_32_0_1_288_2403_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2421:146
  wire [31:0] _delay_fixed_32_0_1_11_2402_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2420:142
  wire [31:0] _delay_fixed_32_0_1_1149_2401_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2419:150
  wire [31:0] _delay_fixed_32_0_1_1291_2400_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2418:150
  wire [31:0] _delay_fixed_32_0_1_11_2399_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2417:142
  wire [31:0] _delay_fixed_32_0_1_1120_2398_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2416:150
  wire [31:0] _delay_fixed_32_0_1_1293_2397_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2415:150
  wire [31:0] _delay_fixed_32_0_1_48_2396_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2414:142
  wire [31:0] _delay_fixed_32_0_1_1261_2395_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2413:150
  wire [31:0] _delay_fixed_32_0_1_1357_2394_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2412:150
  wire [31:0] _delay_fixed_32_0_1_96_2393_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2411:142
  wire [31:0] _delay_fixed_32_0_1_1227_2392_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2410:150
  wire [31:0] _delay_fixed_32_0_1_1410_2391_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2409:150
  wire        _delay_fixed_1_0_0_101_2390_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2408:142
  wire [31:0] _delay_fixed_32_0_1_59_2389_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2407:142
  wire [31:0] _delay_fixed_32_0_1_1496_2388_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2406:150
  wire [31:0] _delay_fixed_32_0_1_1551_2387_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2405:150
  wire [31:0] _delay_fixed_32_0_1_55_2386_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2404:142
  wire [31:0] _delay_fixed_32_0_1_1462_2385_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2403:150
  wire [31:0] _delay_fixed_32_0_1_1602_2384_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2402:150
  wire        _delay_fixed_1_0_0_101_2383_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2401:142
  wire [31:0] _delay_fixed_32_0_1_18_2382_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2400:142
  wire [31:0] _delay_fixed_32_0_1_1463_2381_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2399:150
  wire [31:0] _delay_fixed_32_0_1_1519_2380_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2398:150
  wire [31:0] _delay_fixed_32_0_1_56_2379_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2397:142
  wire [31:0] _delay_fixed_32_0_1_1429_2378_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2396:150
  wire [31:0] _delay_fixed_32_0_1_1540_2377_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2395:150
  wire        _delay_fixed_1_0_0_64_2376_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2394:138
  wire [31:0] _delay_fixed_32_0_1_159_2375_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2393:146
  wire [31:0] _delay_fixed_32_0_1_1360_2374_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2392:150
  wire [31:0] _delay_fixed_32_0_1_1391_2373_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2391:150
  wire [31:0] _delay_fixed_32_0_1_31_2372_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2390:142
  wire [31:0] _delay_fixed_32_0_1_1326_2371_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2389:150
  wire [31:0] _delay_fixed_32_0_1_1450_2370_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2388:150
  wire        _delay_fixed_1_0_0_114_2369_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2387:142
  wire [31:0] _delay_fixed_32_0_1_159_2368_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2386:146
  wire [31:0] _delay_fixed_32_0_1_1394_2367_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2385:150
  wire [31:0] _delay_fixed_32_0_1_1449_2366_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2384:150
  wire [31:0] _delay_fixed_32_0_1_55_2365_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2383:142
  wire [31:0] _delay_fixed_32_0_1_1360_2364_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2382:150
  wire [31:0] _delay_fixed_32_0_1_1487_2363_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2381:150
  wire        _delay_fixed_1_0_0_71_2362_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2380:138
  wire [31:0] _delay_fixed_32_0_1_18_2361_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2379:142
  wire [31:0] _delay_fixed_32_0_1_1520_2360_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2378:150
  wire [31:0] _delay_fixed_32_0_1_1555_2359_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2377:150
  wire [31:0] _delay_fixed_32_0_1_35_2358_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2376:142
  wire [31:0] _delay_fixed_32_0_1_1486_2357_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2375:150
  wire [31:0] _delay_fixed_32_0_1_1604_2356_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2374:150
  wire        _delay_fixed_1_0_0_48_2355_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2373:138
  wire [31:0] _delay_fixed_32_0_1_59_2354_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2372:142
  wire [31:0] _delay_fixed_32_0_1_1557_2353_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2371:150
  wire [31:0] _delay_fixed_32_0_1_1602_2352_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2370:150
  wire [31:0] _delay_fixed_32_0_1_45_2351_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2369:142
  wire [31:0] _delay_fixed_32_0_1_1523_2350_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2368:150
  wire [31:0] _delay_fixed_32_0_1_1626_2349_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2367:150
  wire        _delay_fixed_1_0_0_43_2348_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2366:138
  wire [31:0] _delay_fixed_32_0_1_48_2347_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2365:142
  wire [31:0] _delay_fixed_32_0_1_1268_2346_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2364:150
  wire [31:0] _delay_fixed_32_0_1_1320_2345_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2363:150
  wire [31:0] _delay_fixed_32_0_1_52_2344_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2362:142
  wire [31:0] _delay_fixed_32_0_1_1234_2343_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2361:150
  wire [31:0] _delay_fixed_32_0_1_1306_2342_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2360:150
  wire        _delay_fixed_1_0_0_55_2341_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2359:138
  wire [31:0] _delay_fixed_32_0_1_902_2340_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2358:146
  wire [31:0] _delay_fixed_32_0_1_13_2339_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2357:142
  wire [31:0] _delay_fixed_32_0_1_772_2338_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2356:146
  wire [31:0] _delay_fixed_32_0_1_778_2337_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2355:146
  wire [31:0] _delay_fixed_32_0_1_708_2336_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2354:146
  wire [31:0] _delay_fixed_32_0_1_152_2335_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2353:146
  wire [31:0] _delay_fixed_32_0_1_765_2334_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2352:146
  wire [31:0] _delay_fixed_32_0_1_163_2333_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2351:146
  wire [31:0] _delay_fixed_32_0_1_45_2332_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2350:142
  wire [31:0] _delay_fixed_32_0_1_779_2331_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2349:146
  wire [31:0] _delay_fixed_32_0_1_666_2330_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2348:146
  wire [31:0] _delay_fixed_32_0_1_668_2329_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2347:146
  wire [31:0] _delay_fixed_32_0_1_92_2328_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2346:142
  wire [31:0] _delay_fixed_32_0_1_681_2327_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2345:146
  wire [31:0] _delay_fixed_32_0_1_171_2326_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2344:146
  wire [31:0] _delay_fixed_32_0_1_160_2325_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2343:146
  wire [31:0] _delay_fixed_32_0_1_160_2324_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2342:146
  wire [31:0] _delay_fixed_32_0_1_153_2323_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2341:146
  wire [31:0] _delay_fixed_32_0_1_825_2322_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2340:146
  wire [31:0] _delay_fixed_32_0_1_732_2321_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2339:146
  wire [31:0] _delay_fixed_32_0_1_644_2320_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2338:146
  wire [31:0] _delay_fixed_32_0_1_274_2319_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2337:146
  wire [31:0] _delay_fixed_32_0_1_853_2318_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2336:146
  wire [31:0] _delay_fixed_32_0_1_109_2317_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2335:146
  wire [31:0] _delay_fixed_32_0_1_11_2316_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2334:142
  wire [31:0] _delay_fixed_32_0_1_11_2315_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2333:142
  wire [31:0] _delay_fixed_32_0_1_27_2314_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2332:142
  wire [31:0] _delay_fixed_32_0_1_27_2313_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2331:142
  wire [31:0] _delay_fixed_32_0_1_119_2312_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2330:146
  wire [31:0] _delay_fixed_32_0_1_119_2311_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2329:146
  wire [31:0] _delay_fixed_32_0_1_49_2310_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2328:142
  wire [31:0] _delay_fixed_32_0_1_49_2309_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2327:142
  wire [31:0] _delay_fixed_32_0_1_172_2308_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2326:146
  wire [31:0] _delay_fixed_32_0_1_1316_2307_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2325:150
  wire [31:0] _delay_fixed_32_0_1_1391_2306_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2324:150
  wire [31:0] _delay_fixed_32_0_1_172_2305_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2323:146
  wire [31:0] _delay_fixed_32_0_1_1323_2304_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2322:150
  wire [31:0] _delay_fixed_32_0_1_1488_2303_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2321:150
  wire [31:0] _delay_fixed_32_0_1_6_2302_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2320:138
  wire [31:0] _delay_fixed_32_0_1_1301_2301_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2319:150
  wire [31:0] _delay_fixed_32_0_1_1354_2300_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2318:150
  wire [31:0] _delay_fixed_32_0_1_53_2299_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2317:142
  wire [31:0] _delay_fixed_32_0_1_1267_2298_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2316:150
  wire [31:0] _delay_fixed_32_0_1_1341_2297_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2315:150
  wire        _delay_fixed_1_0_0_63_2296_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2314:138
  wire [31:0] _delay_fixed_32_0_1_248_2295_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2313:146
  wire [31:0] _delay_fixed_32_0_1_1643_2294_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2312:150
  wire [31:0] _delay_fixed_32_0_1_23_2293_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2311:142
  wire [31:0] _delay_fixed_32_0_1_1402_2292_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2310:150
  wire [31:0] _delay_fixed_32_0_1_1408_2291_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2309:150
  wire [31:0] _delay_fixed_32_0_1_6_2290_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2308:138
  wire [31:0] _delay_fixed_32_0_1_1368_2289_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2307:150
  wire [31:0] _delay_fixed_32_0_1_1449_2288_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2306:150
  wire [31:0] _delay_fixed_32_0_1_26_2287_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2305:142
  wire [31:0] _delay_fixed_32_0_1_1662_2286_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2304:150
  wire [31:0] _delay_fixed_32_0_1_1675_2285_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2303:150
  wire [31:0] _delay_fixed_32_0_1_13_2284_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2302:142
  wire [31:0] _delay_fixed_32_0_1_1628_2283_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2301:150
  wire [31:0] _delay_fixed_32_0_1_1691_2282_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2300:150
  wire        _delay_fixed_1_0_0_25_2281_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2299:138
  wire [31:0] _delay_fixed_32_0_1_248_2280_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2298:146
  wire [31:0] _delay_fixed_32_0_1_1666_2279_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2297:150
  wire [31:0] _delay_fixed_32_0_1_1741_2278_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2296:150
  wire [31:0] _delay_fixed_32_0_1_75_2277_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2295:142
  wire [31:0] _delay_fixed_32_0_1_1632_2276_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2294:150
  wire [31:0] _delay_fixed_32_0_1_1771_2275_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2293:150
  wire        _delay_fixed_1_0_0_114_2274_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2292:142
  wire [31:0] _delay_fixed_32_0_1_6_2273_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2291:138
  wire [31:0] _delay_fixed_32_0_1_1338_2272_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2290:150
  wire [31:0] _delay_fixed_32_0_1_1369_2271_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2289:150
  wire [31:0] _delay_fixed_32_0_1_31_2270_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2288:142
  wire [31:0] _delay_fixed_32_0_1_1304_2269_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2287:150
  wire [31:0] _delay_fixed_32_0_1_1392_2268_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2286:150
  wire        _delay_fixed_1_0_0_42_2267_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2285:138
  wire [31:0] _delay_fixed_32_0_1_923_2266_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2284:146
  wire [31:0] _delay_fixed_32_0_1_32_2265_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2283:142
  wire [31:0] _delay_fixed_32_0_1_886_2264_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2282:146
  wire [31:0] _delay_fixed_32_0_1_838_2263_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2281:146
  wire [31:0] _delay_fixed_32_0_1_837_2262_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2280:146
  wire [31:0] _delay_fixed_32_0_1_155_2261_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2279:146
  wire [31:0] _delay_fixed_32_0_1_913_2260_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2278:146
  wire [31:0] _delay_fixed_32_0_1_130_2259_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2277:146
  wire [31:0] _delay_fixed_32_0_1_29_2258_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2276:142
  wire [31:0] _delay_fixed_32_0_1_965_2257_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2275:146
  wire [31:0] _delay_fixed_32_0_1_908_2256_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2274:146
  wire [31:0] _delay_fixed_32_0_1_819_2255_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2273:146
  wire [31:0] _delay_fixed_32_0_1_67_2254_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2272:142
  wire [31:0] _delay_fixed_32_0_1_906_2253_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2271:146
  wire [31:0] _delay_fixed_32_0_1_71_2252_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2270:142
  wire [31:0] _delay_fixed_32_0_1_7_2251_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2269:138
  wire [31:0] _delay_fixed_32_0_1_7_2250_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2268:138
  wire [31:0] _delay_fixed_32_0_1_86_2249_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2267:142
  wire [31:0] _delay_fixed_32_0_1_986_2248_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2266:146
  wire [31:0] _delay_fixed_32_0_1_898_2247_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2265:146
  wire [31:0] _delay_fixed_32_0_1_871_2246_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2264:146
  wire [31:0] _delay_fixed_32_0_1_114_2245_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2263:146
  wire [31:0] _delay_fixed_32_0_1_1013_2244_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2262:150
  wire [31:0] _delay_fixed_32_0_1_17_2243_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2261:142
  wire [31:0] _delay_fixed_32_0_1_145_2242_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2260:146
  wire [31:0] _delay_fixed_32_0_1_145_2241_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2259:146
  wire [31:0] _delay_fixed_32_0_1_71_2240_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2258:142
  wire [31:0] _delay_fixed_32_0_1_71_2239_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2257:142
  wire [31:0] _delay_fixed_32_0_1_65_2238_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2256:142
  wire [31:0] _delay_fixed_32_0_1_65_2237_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2255:142
  wire [31:0] _delay_fixed_32_0_1_102_2236_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2254:146
  wire [31:0] _delay_fixed_32_0_1_102_2235_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2253:146
  wire [31:0] _delay_fixed_32_0_1_21_2234_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2252:142
  wire [31:0] _delay_fixed_32_0_1_1365_2233_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2251:150
  wire [31:0] _delay_fixed_32_0_1_1478_2232_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2250:150
  wire [31:0] _delay_fixed_32_0_1_21_2231_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2249:142
  wire [31:0] _delay_fixed_32_0_1_1421_2230_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2248:150
  wire [31:0] _delay_fixed_32_0_1_1561_2229_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2247:150
  wire [31:0] _delay_fixed_32_0_1_52_2228_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2246:142
  wire [31:0] _delay_fixed_32_0_1_1517_2227_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2245:150
  wire [31:0] _delay_fixed_32_0_1_1579_2226_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2244:150
  wire [31:0] _delay_fixed_32_0_1_62_2225_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2243:142
  wire [31:0] _delay_fixed_32_0_1_1483_2224_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2242:150
  wire [31:0] _delay_fixed_32_0_1_1612_2223_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2241:150
  wire        _delay_fixed_1_0_0_92_2222_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2240:138
  wire [31:0] _delay_fixed_32_0_1_373_2221_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2239:146
  wire [31:0] _delay_fixed_32_0_1_1756_2220_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2238:150
  wire [31:0] _delay_fixed_32_0_1_1775_2219_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2237:150
  wire [31:0] _delay_fixed_32_0_1_19_2218_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2236:142
  wire [31:0] _delay_fixed_32_0_1_1722_2217_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2235:150
  wire [31:0] _delay_fixed_32_0_1_1790_2216_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2234:150
  wire        _delay_fixed_1_0_0_5_2215_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2233:134
  wire [31:0] _delay_fixed_32_0_1_388_2214_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2232:146
  wire [31:0] _delay_fixed_32_0_1_1763_2213_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2231:150
  wire [31:0] _delay_fixed_32_0_1_1804_2212_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2230:150
  wire [31:0] _delay_fixed_32_0_1_41_2211_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2229:142
  wire [31:0] _delay_fixed_32_0_1_1729_2210_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2228:150
  wire [31:0] _delay_fixed_32_0_1_1848_2209_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2227:150
  wire        _delay_fixed_1_0_0_86_2208_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2226:138
  wire [31:0] _delay_fixed_32_0_1_84_2207_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2225:142
  wire [31:0] _delay_fixed_32_0_1_1441_2206_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2224:150
  wire [31:0] _delay_fixed_32_0_1_1452_2205_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2223:150
  wire [31:0] _delay_fixed_32_0_1_11_2204_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2222:142
  wire [31:0] _delay_fixed_32_0_1_1407_2203_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2221:150
  wire [31:0] _delay_fixed_32_0_1_1446_2202_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2220:150
  wire [31:0] _delay_fixed_32_0_1_26_2201_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2219:142
  wire [31:0] _delay_fixed_32_0_1_84_2200_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2218:142
  wire [31:0] _delay_fixed_32_0_1_1371_2199_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2217:150
  wire [31:0] _delay_fixed_32_0_1_1391_2198_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2216:150
  wire [31:0] _delay_fixed_32_0_1_20_2197_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2215:142
  wire [31:0] _delay_fixed_32_0_1_1337_2196_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2214:150
  wire [31:0] _delay_fixed_32_0_1_1391_2195_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2213:150
  wire [31:0] _delay_fixed_32_0_1_29_2194_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2212:142
  wire [31:0] _delay_fixed_32_0_1_388_2193_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2211:146
  wire [31:0] _delay_fixed_32_0_1_1865_2192_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2210:150
  wire [31:0] _delay_fixed_32_0_1_1940_2191_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2209:150
  wire [31:0] _delay_fixed_32_0_1_75_2190_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2208:142
  wire [31:0] _delay_fixed_32_0_1_1831_2189_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2207:150
  wire [31:0] _delay_fixed_32_0_1_1996_2188_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2206:150
  wire        _delay_fixed_1_0_0_106_2187_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2205:142
  wire [31:0] _delay_fixed_32_0_1_373_2186_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2204:146
  wire [31:0] _delay_fixed_32_0_1_1719_2185_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2203:150
  wire [31:0] _delay_fixed_32_0_1_1779_2184_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2202:150
  wire [31:0] _delay_fixed_32_0_1_60_2183_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2201:142
  wire [31:0] _delay_fixed_32_0_1_1685_2182_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2200:150
  wire [31:0] _delay_fixed_32_0_1_1812_2181_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2199:150
  wire        _delay_fixed_1_0_0_60_2180_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2198:138
  wire [31:0] _delay_fixed_32_0_1_52_2179_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2197:142
  wire [31:0] _delay_fixed_32_0_1_1535_2178_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2196:150
  wire [31:0] _delay_fixed_32_0_1_1548_2177_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2195:150
  wire [31:0] _delay_fixed_32_0_1_13_2176_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2194:142
  wire [31:0] _delay_fixed_32_0_1_1501_2175_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2193:150
  wire [31:0] _delay_fixed_32_0_1_1596_2174_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2192:150
  wire        _delay_fixed_1_0_0_29_2173_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2191:138
  wire [31:0] _delay_fixed_32_0_1_990_2172_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2190:146
  wire [31:0] _delay_fixed_32_0_1_274_2171_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2189:146
  wire [31:0] _delay_fixed_32_0_1_1154_2170_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2188:150
  wire [31:0] _delay_fixed_32_0_1_1099_2169_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2187:150
  wire [31:0] _delay_fixed_32_0_1_1055_2168_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2186:150
  wire [31:0] _delay_fixed_32_0_1_194_2167_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2185:146
  wire [31:0] _delay_fixed_32_0_1_825_2166_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2184:146
  wire [31:0] _delay_fixed_32_0_1_436_2165_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2183:146
  wire [31:0] _delay_fixed_32_0_1_46_2164_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2182:142
  wire [31:0] _delay_fixed_32_0_1_1041_2163_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2181:150
  wire [31:0] _delay_fixed_32_0_1_1007_2162_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2180:150
  wire [31:0] _delay_fixed_32_0_1_876_2161_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2179:146
  wire [31:0] _delay_fixed_32_0_1_240_2160_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2178:146
  wire [31:0] _delay_fixed_32_0_1_980_2159_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2177:146
  wire [31:0] _delay_fixed_32_0_1_147_2158_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2176:146
  wire [31:0] _delay_fixed_32_0_1_16_2157_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2175:142
  wire [31:0] _delay_fixed_32_0_1_16_2156_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2174:142
  wire [31:0] _delay_fixed_32_0_1_156_2155_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2173:146
  wire [31:0] _delay_fixed_32_0_1_962_2154_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2172:146
  wire [31:0] _delay_fixed_32_0_1_917_2153_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2171:146
  wire [31:0] _delay_fixed_32_0_1_784_2152_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2170:146
  wire [31:0] _delay_fixed_32_0_1_273_2151_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2169:146
  wire [31:0] _delay_fixed_32_0_1_996_2150_out;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2168:146
  wire [31:0] _const2149_const_fix_32_0_1__0000000000000235;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2167:90
  wire [31:0] _const2146_const_fix_32_0_1__00000000000000ff;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2166:90
  wire [31:0] _const2144_const_fix_32_0_1__0000000000000004;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2165:90
  wire [31:0] _const2111_const_fix_32_0_1__0000000000000454;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2164:90
  wire [31:0] _const2106_const_fix_32_0_1__0000000000000080;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2163:90
  wire [31:0] _const2102_const_fix_32_0_1__00000000000000b5;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2162:90
  wire [31:0] _const2098_const_fix_32_0_1__0000000000000ec8;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2161:90
  wire [31:0] _const2097_const_fix_32_0_1__0000000000000968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2160:90
  wire [31:0] _const2086_const_fix_32_0_1__ffffffffffffff00;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2159:90
  wire [31:0] _const2081_const_fix_32_0_1__0000000000000d4e;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2158:90
  wire [31:0] _const2074_const_fix_32_0_1__00000000000008e4;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2157:90
  wire [31:0] _const2068_const_fix_32_0_1__0000000000000fb1;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2156:90
  wire [31:0] _const2065_const_fix_32_0_1__000000000000031f;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2155:90
  wire [31:0] _const2060_const_fix_32_0_1__0000000000000620;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2154:90
  wire [31:0] _const2045_const_fix_32_0_1__0000000000002000;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2153:90
  wire [31:0] _MUX2005__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2151:169
  wire        _LT2004__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2150:139
  wire [31:0] _MUX2003__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2149:169
  wire        _GT2002__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2148:139
  wire [31:0] _dup2001__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2147:154
  wire [31:0] _dup2001__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2147:154
  wire [31:0] _dup2001__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2147:154
  wire [31:0] _SHR142000__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2146:97
  wire [31:0] _SUB1999__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2145:114
  wire [31:0] _MUX1997__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2143:169
  wire        _LT1996__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2142:139
  wire [31:0] _MUX1995__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2141:169
  wire        _GT1994__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2140:139
  wire [31:0] _dup1993__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2139:154
  wire [31:0] _dup1993__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2139:154
  wire [31:0] _dup1993__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2139:154
  wire [31:0] _SHR141992__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2138:97
  wire [31:0] _SUB1991__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2137:114
  wire [31:0] _MUX1989__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2135:169
  wire        _LT1988__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2134:139
  wire [31:0] _MUX1987__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2133:169
  wire        _GT1986__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2132:139
  wire [31:0] _dup1985__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2131:154
  wire [31:0] _dup1985__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2131:154
  wire [31:0] _dup1985__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2131:154
  wire [31:0] _SHR141984__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2130:97
  wire [31:0] _SUB1983__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2129:114
  wire [31:0] _MUX1981__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2127:169
  wire        _LT1980__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2126:139
  wire [31:0] _MUX1979__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2125:169
  wire        _GT1978__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2124:139
  wire [31:0] _dup1977__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2123:154
  wire [31:0] _dup1977__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2123:154
  wire [31:0] _dup1977__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2123:154
  wire [31:0] _SHR141976__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2122:97
  wire [31:0] _SUB1975__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2121:114
  wire [31:0] _MUX1973__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2119:169
  wire        _LT1972__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2118:139
  wire [31:0] _MUX1971__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2117:169
  wire        _GT1970__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2116:139
  wire [31:0] _dup1969__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2115:154
  wire [31:0] _dup1969__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2115:154
  wire [31:0] _dup1969__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2115:154
  wire [31:0] _SHR141968__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2114:97
  wire [31:0] _ADD1967__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2113:135
  wire [31:0] _dup1966__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2112:116
  wire [31:0] _dup1966__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2112:116
  wire [31:0] _dup1965__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2111:116
  wire [31:0] _dup1965__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2111:116
  wire [31:0] _MUX1963__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2109:169
  wire        _LT1962__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2108:139
  wire [31:0] _MUX1961__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2107:169
  wire        _GT1960__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2106:139
  wire [31:0] _dup1959__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2105:154
  wire [31:0] _dup1959__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2105:154
  wire [31:0] _dup1959__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2105:154
  wire [31:0] _SHR141958__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2104:97
  wire [31:0] _ADD1957__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2103:135
  wire [31:0] _dup1956__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2102:116
  wire [31:0] _dup1956__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2102:116
  wire [31:0] _dup1955__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2101:116
  wire [31:0] _dup1955__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2101:116
  wire [31:0] _MUX1953__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2099:169
  wire        _LT1952__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2098:139
  wire [31:0] _MUX1951__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2097:169
  wire        _GT1950__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2096:139
  wire [31:0] _dup1949__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2095:154
  wire [31:0] _dup1949__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2095:154
  wire [31:0] _dup1949__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2095:154
  wire [31:0] _SHR141948__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2094:97
  wire [31:0] _ADD1947__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2093:135
  wire [31:0] _dup1946__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2092:116
  wire [31:0] _dup1946__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2092:116
  wire [31:0] _dup1945__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2091:116
  wire [31:0] _dup1945__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2091:116
  wire [31:0] _MUX1943__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2089:169
  wire        _LT1942__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2088:139
  wire [31:0] _MUX1941__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2087:169
  wire        _GT1940__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2086:139
  wire [31:0] _dup1939__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2085:154
  wire [31:0] _dup1939__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2085:154
  wire [31:0] _dup1939__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2085:154
  wire [31:0] _SHR141938__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2084:97
  wire [31:0] _ADD1937__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2083:135
  wire [31:0] _dup1936__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2082:116
  wire [31:0] _dup1936__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2082:116
  wire [31:0] _dup1935__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2081:116
  wire [31:0] _dup1935__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2081:116
  wire [31:0] _SHR81934__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2080:91
  wire [31:0] _ADD1933__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2079:135
  wire [31:0] _MUL1932__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2078:136
  wire [31:0] _SUB1931__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2077:114
  wire [31:0] _SHR81930__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2076:91
  wire [31:0] _ADD1929__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2075:135
  wire [31:0] _MUL1928__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2074:136
  wire [31:0] _ADD1927__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2073:135
  wire [31:0] _dup1926__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2072:116
  wire [31:0] _dup1926__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2072:116
  wire [31:0] _dup1925__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2071:116
  wire [31:0] _dup1925__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2071:116
  wire [31:0] _SUB1924__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2070:114
  wire [31:0] _ADD1923__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2069:135
  wire [31:0] _dup1922__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2068:116
  wire [31:0] _dup1922__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2068:116
  wire [31:0] _dup1921__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2067:116
  wire [31:0] _dup1921__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2067:116
  wire [31:0] _SUB1920__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2066:114
  wire [31:0] _ADD1919__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2065:135
  wire [31:0] _dup1918__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2064:116
  wire [31:0] _dup1918__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2064:116
  wire [31:0] _dup1917__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2063:116
  wire [31:0] _dup1917__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2063:116
  wire [31:0] _SUB1916__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2062:114
  wire [31:0] _ADD1915__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2061:135
  wire [31:0] _dup1914__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2060:116
  wire [31:0] _dup1914__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2060:116
  wire [31:0] _dup1913__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2059:116
  wire [31:0] _dup1913__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2059:116
  wire [31:0] _SUB1912__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2058:114
  wire [31:0] _ADD1911__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2057:135
  wire [31:0] _dup1910__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2056:116
  wire [31:0] _dup1910__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2056:116
  wire [31:0] _dup1909__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2055:116
  wire [31:0] _dup1909__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2055:116
  wire [31:0] _SHR31908__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2054:93
  wire [31:0] _ADD1907__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2053:135
  wire [31:0] _MUL1906__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2052:136
  wire [31:0] _SHR31905__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2051:93
  wire [31:0] _SUB1904__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2050:114
  wire [31:0] _dup1903__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2049:116
  wire [31:0] _dup1903__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2049:116
  wire [31:0] _MUL1902__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2048:136
  wire [31:0] _ADD1901__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2047:135
  wire [31:0] _MUL1900__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2046:136
  wire [31:0] _ADD1899__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2045:135
  wire [31:0] _dup1898__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2044:116
  wire [31:0] _dup1898__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2044:116
  wire [31:0] _dup1897__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2043:116
  wire [31:0] _dup1897__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2043:116
  wire [31:0] _SUB1896__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2042:114
  wire [31:0] _ADD1895__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2041:135
  wire [31:0] _dup1894__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2040:116
  wire [31:0] _dup1894__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2040:116
  wire [31:0] _dup1893__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2039:116
  wire [31:0] _dup1893__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2039:116
  wire [31:0] _SHR31892__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2038:93
  wire [31:0] _SUB1891__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2037:114
  wire [31:0] _MUL1890__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2036:136
  wire [31:0] _SHR31889__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2035:93
  wire [31:0] _SUB1888__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2034:114
  wire [31:0] _dup1887__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2033:116
  wire [31:0] _dup1887__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2033:116
  wire [31:0] _MUL1886__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2032:136
  wire [31:0] _ADD1885__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2031:135
  wire [31:0] _MUL1884__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2030:136
  wire [31:0] _ADD1883__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2029:135
  wire [31:0] _dup1882__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2028:116
  wire [31:0] _dup1882__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2028:116
  wire [31:0] _dup1881__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2027:116
  wire [31:0] _dup1881__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2027:116
  wire [31:0] _SHR31880__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2026:93
  wire [31:0] _SUB1879__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2025:114
  wire [31:0] _MUL1878__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2024:136
  wire [31:0] _SHR31877__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2023:93
  wire [31:0] _ADD1876__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2022:135
  wire [31:0] _dup1875__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2021:116
  wire [31:0] _dup1875__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2021:116
  wire [31:0] _MUL1874__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2020:136
  wire [31:0] _ADD1873__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2019:135
  wire [31:0] _MUL1872__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2018:136
  wire [31:0] _ADD1871__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2017:135
  wire [31:0] _dup1870__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2016:116
  wire [31:0] _dup1870__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2016:116
  wire [31:0] _dup1869__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2015:116
  wire [31:0] _dup1869__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2015:116
  wire [31:0] _ADD1868__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2014:135
  wire [31:0] _SHL81867__dfc_wire_1923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2013:93
  wire [31:0] _CAST1866__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2012:88
  wire [31:0] _CAST1865__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2011:88
  wire [31:0] _CAST1864__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2010:88
  wire [31:0] _CAST1863__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2009:88
  wire [31:0] _CAST1862__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2008:88
  wire [31:0] _CAST1861__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2007:88
  wire [31:0] _CAST1860__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2006:88
  wire [31:0] _SHL81859__dfc_wire_1923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2005:93
  wire [31:0] _CAST1858__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2004:88
  wire [31:0] _MUX1856__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2002:169
  wire        _LT1855__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2001:139
  wire [31:0] _MUX1854__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2000:169
  wire        _GT1853__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1999:139
  wire [31:0] _dup1852__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1998:154
  wire [31:0] _dup1852__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1998:154
  wire [31:0] _dup1852__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1998:154
  wire [31:0] _SHR141851__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1997:97
  wire [31:0] _SUB1850__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1996:114
  wire [31:0] _MUX1848__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1994:169
  wire        _LT1847__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1993:139
  wire [31:0] _MUX1846__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1992:169
  wire        _GT1845__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1991:139
  wire [31:0] _dup1844__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1990:154
  wire [31:0] _dup1844__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1990:154
  wire [31:0] _dup1844__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1990:154
  wire [31:0] _SHR141843__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1989:97
  wire [31:0] _SUB1842__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1988:114
  wire [31:0] _MUX1840__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1986:169
  wire        _LT1839__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1985:139
  wire [31:0] _MUX1838__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1984:169
  wire        _GT1837__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1983:139
  wire [31:0] _dup1836__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1982:154
  wire [31:0] _dup1836__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1982:154
  wire [31:0] _dup1836__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1982:154
  wire [31:0] _SHR141835__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1981:97
  wire [31:0] _SUB1834__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1980:114
  wire [31:0] _MUX1832__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1978:169
  wire        _LT1831__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1977:139
  wire [31:0] _MUX1830__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1976:169
  wire        _GT1829__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1975:139
  wire [31:0] _dup1828__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1974:154
  wire [31:0] _dup1828__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1974:154
  wire [31:0] _dup1828__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1974:154
  wire [31:0] _SHR141827__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1973:97
  wire [31:0] _SUB1826__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1972:114
  wire [31:0] _MUX1824__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1970:169
  wire        _LT1823__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1969:139
  wire [31:0] _MUX1822__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1968:169
  wire        _GT1821__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1967:139
  wire [31:0] _dup1820__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1966:154
  wire [31:0] _dup1820__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1966:154
  wire [31:0] _dup1820__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1966:154
  wire [31:0] _SHR141819__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1965:97
  wire [31:0] _ADD1818__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1964:135
  wire [31:0] _dup1817__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1963:116
  wire [31:0] _dup1817__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1963:116
  wire [31:0] _dup1816__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1962:116
  wire [31:0] _dup1816__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1962:116
  wire [31:0] _MUX1814__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1960:169
  wire        _LT1813__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1959:139
  wire [31:0] _MUX1812__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1958:169
  wire        _GT1811__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1957:139
  wire [31:0] _dup1810__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1956:154
  wire [31:0] _dup1810__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1956:154
  wire [31:0] _dup1810__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1956:154
  wire [31:0] _SHR141809__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1955:97
  wire [31:0] _ADD1808__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1954:135
  wire [31:0] _dup1807__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1953:116
  wire [31:0] _dup1807__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1953:116
  wire [31:0] _dup1806__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1952:116
  wire [31:0] _dup1806__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1952:116
  wire [31:0] _MUX1804__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1950:169
  wire        _LT1803__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1949:139
  wire [31:0] _MUX1802__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1948:169
  wire        _GT1801__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1947:139
  wire [31:0] _dup1800__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1946:154
  wire [31:0] _dup1800__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1946:154
  wire [31:0] _dup1800__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1946:154
  wire [31:0] _SHR141799__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1945:97
  wire [31:0] _ADD1798__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1944:135
  wire [31:0] _dup1797__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1943:116
  wire [31:0] _dup1797__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1943:116
  wire [31:0] _dup1796__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1942:116
  wire [31:0] _dup1796__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1942:116
  wire [31:0] _MUX1794__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1940:169
  wire        _LT1793__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1939:139
  wire [31:0] _MUX1792__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1938:169
  wire        _GT1791__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1937:139
  wire [31:0] _dup1790__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1936:154
  wire [31:0] _dup1790__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1936:154
  wire [31:0] _dup1790__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1936:154
  wire [31:0] _SHR141789__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1935:97
  wire [31:0] _ADD1788__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1934:135
  wire [31:0] _dup1787__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1933:116
  wire [31:0] _dup1787__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1933:116
  wire [31:0] _dup1786__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1932:116
  wire [31:0] _dup1786__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1932:116
  wire [31:0] _SHR81785__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1931:91
  wire [31:0] _ADD1784__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1930:135
  wire [31:0] _MUL1783__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1929:136
  wire [31:0] _SUB1782__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1928:114
  wire [31:0] _SHR81781__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1927:91
  wire [31:0] _ADD1780__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1926:135
  wire [31:0] _MUL1779__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1925:136
  wire [31:0] _ADD1778__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1924:135
  wire [31:0] _dup1777__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1923:116
  wire [31:0] _dup1777__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1923:116
  wire [31:0] _dup1776__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1922:116
  wire [31:0] _dup1776__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1922:116
  wire [31:0] _SUB1775__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1921:114
  wire [31:0] _ADD1774__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1920:135
  wire [31:0] _dup1773__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1919:116
  wire [31:0] _dup1773__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1919:116
  wire [31:0] _dup1772__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1918:116
  wire [31:0] _dup1772__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1918:116
  wire [31:0] _SUB1771__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1917:114
  wire [31:0] _ADD1770__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1916:135
  wire [31:0] _dup1769__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1915:116
  wire [31:0] _dup1769__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1915:116
  wire [31:0] _dup1768__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1914:116
  wire [31:0] _dup1768__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1914:116
  wire [31:0] _SUB1767__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1913:114
  wire [31:0] _ADD1766__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1912:135
  wire [31:0] _dup1765__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1911:116
  wire [31:0] _dup1765__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1911:116
  wire [31:0] _dup1764__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1910:116
  wire [31:0] _dup1764__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1910:116
  wire [31:0] _SUB1763__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1909:114
  wire [31:0] _ADD1762__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1908:135
  wire [31:0] _dup1761__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1907:116
  wire [31:0] _dup1761__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1907:116
  wire [31:0] _dup1760__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1906:116
  wire [31:0] _dup1760__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1906:116
  wire [31:0] _SHR31759__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1905:93
  wire [31:0] _ADD1758__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1904:135
  wire [31:0] _MUL1757__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1903:136
  wire [31:0] _SHR31756__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1902:93
  wire [31:0] _SUB1755__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1901:114
  wire [31:0] _dup1754__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1900:116
  wire [31:0] _dup1754__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1900:116
  wire [31:0] _MUL1753__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1899:136
  wire [31:0] _ADD1752__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1898:135
  wire [31:0] _MUL1751__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1897:136
  wire [31:0] _ADD1750__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1896:135
  wire [31:0] _dup1749__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1895:116
  wire [31:0] _dup1749__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1895:116
  wire [31:0] _dup1748__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1894:116
  wire [31:0] _dup1748__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1894:116
  wire [31:0] _SUB1747__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1893:114
  wire [31:0] _ADD1746__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1892:135
  wire [31:0] _dup1745__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1891:116
  wire [31:0] _dup1745__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1891:116
  wire [31:0] _dup1744__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1890:116
  wire [31:0] _dup1744__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1890:116
  wire [31:0] _SHR31743__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1889:93
  wire [31:0] _SUB1742__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1888:114
  wire [31:0] _MUL1741__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1887:136
  wire [31:0] _SHR31740__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1886:93
  wire [31:0] _SUB1739__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1885:114
  wire [31:0] _dup1738__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1884:116
  wire [31:0] _dup1738__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1884:116
  wire [31:0] _MUL1737__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1883:136
  wire [31:0] _ADD1736__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1882:135
  wire [31:0] _MUL1735__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1881:136
  wire [31:0] _ADD1734__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1880:135
  wire [31:0] _dup1733__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1879:116
  wire [31:0] _dup1733__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1879:116
  wire [31:0] _dup1732__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1878:116
  wire [31:0] _dup1732__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1878:116
  wire [31:0] _SHR31731__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1877:93
  wire [31:0] _SUB1730__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1876:114
  wire [31:0] _MUL1729__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1875:136
  wire [31:0] _SHR31728__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1874:93
  wire [31:0] _ADD1727__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1873:135
  wire [31:0] _dup1726__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1872:116
  wire [31:0] _dup1726__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1872:116
  wire [31:0] _MUL1725__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1871:136
  wire [31:0] _ADD1724__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1870:135
  wire [31:0] _MUL1723__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1869:136
  wire [31:0] _ADD1722__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1868:135
  wire [31:0] _dup1721__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1867:116
  wire [31:0] _dup1721__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1867:116
  wire [31:0] _dup1720__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1866:116
  wire [31:0] _dup1720__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1866:116
  wire [31:0] _ADD1719__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1865:135
  wire [31:0] _SHL81718__dfc_wire_1923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1864:93
  wire [31:0] _CAST1717__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1863:88
  wire [31:0] _CAST1716__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1862:88
  wire [31:0] _CAST1715__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1861:88
  wire [31:0] _CAST1714__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1860:88
  wire [31:0] _CAST1713__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1859:88
  wire [31:0] _CAST1712__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1858:88
  wire [31:0] _CAST1711__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1857:88
  wire [31:0] _SHL81710__dfc_wire_1923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1856:93
  wire [31:0] _CAST1709__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1855:88
  wire [31:0] _MUX1707__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1853:169
  wire        _LT1706__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1852:139
  wire [31:0] _MUX1705__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1851:169
  wire        _GT1704__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1850:139
  wire [31:0] _dup1703__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1849:154
  wire [31:0] _dup1703__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1849:154
  wire [31:0] _dup1703__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1849:154
  wire [31:0] _SHR141702__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1848:97
  wire [31:0] _SUB1701__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1847:114
  wire [31:0] _MUX1699__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1845:169
  wire        _LT1698__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1844:139
  wire [31:0] _MUX1697__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1843:169
  wire        _GT1696__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1842:139
  wire [31:0] _dup1695__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1841:154
  wire [31:0] _dup1695__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1841:154
  wire [31:0] _dup1695__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1841:154
  wire [31:0] _SHR141694__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1840:97
  wire [31:0] _SUB1693__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1839:114
  wire [31:0] _MUX1691__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1837:169
  wire        _LT1690__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1836:139
  wire [31:0] _MUX1689__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1835:169
  wire        _GT1688__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1834:139
  wire [31:0] _dup1687__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1833:154
  wire [31:0] _dup1687__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1833:154
  wire [31:0] _dup1687__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1833:154
  wire [31:0] _SHR141686__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1832:97
  wire [31:0] _SUB1685__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1831:114
  wire [31:0] _MUX1683__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1829:169
  wire        _LT1682__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1828:139
  wire [31:0] _MUX1681__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1827:169
  wire        _GT1680__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1826:139
  wire [31:0] _dup1679__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1825:154
  wire [31:0] _dup1679__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1825:154
  wire [31:0] _dup1679__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1825:154
  wire [31:0] _SHR141678__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1824:97
  wire [31:0] _SUB1677__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1823:114
  wire [31:0] _MUX1675__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1821:169
  wire        _LT1674__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1820:139
  wire [31:0] _MUX1673__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1819:169
  wire        _GT1672__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1818:139
  wire [31:0] _dup1671__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1817:154
  wire [31:0] _dup1671__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1817:154
  wire [31:0] _dup1671__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1817:154
  wire [31:0] _SHR141670__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1816:97
  wire [31:0] _ADD1669__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1815:135
  wire [31:0] _dup1668__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1814:116
  wire [31:0] _dup1668__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1814:116
  wire [31:0] _dup1667__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1813:116
  wire [31:0] _dup1667__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1813:116
  wire [31:0] _MUX1665__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1811:169
  wire        _LT1664__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1810:139
  wire [31:0] _MUX1663__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1809:169
  wire        _GT1662__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1808:139
  wire [31:0] _dup1661__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1807:154
  wire [31:0] _dup1661__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1807:154
  wire [31:0] _dup1661__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1807:154
  wire [31:0] _SHR141660__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1806:97
  wire [31:0] _ADD1659__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1805:135
  wire [31:0] _dup1658__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1804:116
  wire [31:0] _dup1658__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1804:116
  wire [31:0] _dup1657__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1803:116
  wire [31:0] _dup1657__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1803:116
  wire [31:0] _MUX1655__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1801:169
  wire        _LT1654__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1800:139
  wire [31:0] _MUX1653__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1799:169
  wire        _GT1652__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1798:139
  wire [31:0] _dup1651__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1797:154
  wire [31:0] _dup1651__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1797:154
  wire [31:0] _dup1651__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1797:154
  wire [31:0] _SHR141650__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1796:97
  wire [31:0] _ADD1649__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1795:135
  wire [31:0] _dup1648__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1794:116
  wire [31:0] _dup1648__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1794:116
  wire [31:0] _dup1647__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1793:116
  wire [31:0] _dup1647__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1793:116
  wire [31:0] _MUX1645__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1791:169
  wire        _LT1644__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1790:139
  wire [31:0] _MUX1643__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1789:169
  wire        _GT1642__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1788:139
  wire [31:0] _dup1641__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1787:154
  wire [31:0] _dup1641__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1787:154
  wire [31:0] _dup1641__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1787:154
  wire [31:0] _SHR141640__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1786:97
  wire [31:0] _ADD1639__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1785:135
  wire [31:0] _dup1638__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1784:116
  wire [31:0] _dup1638__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1784:116
  wire [31:0] _dup1637__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1783:116
  wire [31:0] _dup1637__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1783:116
  wire [31:0] _SHR81636__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1782:91
  wire [31:0] _ADD1635__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1781:135
  wire [31:0] _MUL1634__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1780:136
  wire [31:0] _SUB1633__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1779:114
  wire [31:0] _SHR81632__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1778:91
  wire [31:0] _ADD1631__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1777:135
  wire [31:0] _MUL1630__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1776:136
  wire [31:0] _ADD1629__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1775:135
  wire [31:0] _dup1628__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1774:116
  wire [31:0] _dup1628__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1774:116
  wire [31:0] _dup1627__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1773:116
  wire [31:0] _dup1627__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1773:116
  wire [31:0] _SUB1626__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1772:114
  wire [31:0] _ADD1625__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1771:135
  wire [31:0] _dup1624__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1770:116
  wire [31:0] _dup1624__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1770:116
  wire [31:0] _dup1623__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1769:116
  wire [31:0] _dup1623__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1769:116
  wire [31:0] _SUB1622__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1768:114
  wire [31:0] _ADD1621__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1767:135
  wire [31:0] _dup1620__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1766:116
  wire [31:0] _dup1620__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1766:116
  wire [31:0] _dup1619__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1765:116
  wire [31:0] _dup1619__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1765:116
  wire [31:0] _SUB1618__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1764:114
  wire [31:0] _ADD1617__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1763:135
  wire [31:0] _dup1616__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1762:116
  wire [31:0] _dup1616__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1762:116
  wire [31:0] _dup1615__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1761:116
  wire [31:0] _dup1615__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1761:116
  wire [31:0] _SUB1614__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1760:114
  wire [31:0] _ADD1613__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1759:135
  wire [31:0] _dup1612__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1758:116
  wire [31:0] _dup1612__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1758:116
  wire [31:0] _dup1611__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1757:116
  wire [31:0] _dup1611__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1757:116
  wire [31:0] _SHR31610__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1756:93
  wire [31:0] _ADD1609__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1755:135
  wire [31:0] _MUL1608__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1754:136
  wire [31:0] _SHR31607__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1753:93
  wire [31:0] _SUB1606__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1752:114
  wire [31:0] _dup1605__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1751:116
  wire [31:0] _dup1605__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1751:116
  wire [31:0] _MUL1604__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1750:136
  wire [31:0] _ADD1603__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1749:135
  wire [31:0] _MUL1602__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1748:136
  wire [31:0] _ADD1601__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1747:135
  wire [31:0] _dup1600__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1746:116
  wire [31:0] _dup1600__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1746:116
  wire [31:0] _dup1599__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1745:116
  wire [31:0] _dup1599__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1745:116
  wire [31:0] _SUB1598__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1744:114
  wire [31:0] _ADD1597__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1743:135
  wire [31:0] _dup1596__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1742:116
  wire [31:0] _dup1596__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1742:116
  wire [31:0] _dup1595__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1741:116
  wire [31:0] _dup1595__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1741:116
  wire [31:0] _SHR31594__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1740:93
  wire [31:0] _SUB1593__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1739:114
  wire [31:0] _MUL1592__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1738:136
  wire [31:0] _SHR31591__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1737:93
  wire [31:0] _SUB1590__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1736:114
  wire [31:0] _dup1589__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1735:116
  wire [31:0] _dup1589__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1735:116
  wire [31:0] _MUL1588__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1734:136
  wire [31:0] _ADD1587__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1733:135
  wire [31:0] _MUL1586__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1732:136
  wire [31:0] _ADD1585__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1731:135
  wire [31:0] _dup1584__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1730:116
  wire [31:0] _dup1584__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1730:116
  wire [31:0] _dup1583__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1729:116
  wire [31:0] _dup1583__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1729:116
  wire [31:0] _SHR31582__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1728:93
  wire [31:0] _SUB1581__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1727:114
  wire [31:0] _MUL1580__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1726:136
  wire [31:0] _SHR31579__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1725:93
  wire [31:0] _ADD1578__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1724:135
  wire [31:0] _dup1577__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1723:116
  wire [31:0] _dup1577__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1723:116
  wire [31:0] _MUL1576__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1722:136
  wire [31:0] _ADD1575__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1721:135
  wire [31:0] _MUL1574__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1720:136
  wire [31:0] _ADD1573__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1719:135
  wire [31:0] _dup1572__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1718:116
  wire [31:0] _dup1572__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1718:116
  wire [31:0] _dup1571__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1717:116
  wire [31:0] _dup1571__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1717:116
  wire [31:0] _ADD1570__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1716:135
  wire [31:0] _SHL81569__dfc_wire_1923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1715:93
  wire [31:0] _CAST1568__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1714:88
  wire [31:0] _CAST1567__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1713:88
  wire [31:0] _CAST1566__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1712:88
  wire [31:0] _CAST1565__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1711:88
  wire [31:0] _CAST1564__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1710:88
  wire [31:0] _CAST1563__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1709:88
  wire [31:0] _CAST1562__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1708:88
  wire [31:0] _SHL81561__dfc_wire_1923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1707:93
  wire [31:0] _CAST1560__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1706:88
  wire [31:0] _MUX1558__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1704:169
  wire        _LT1557__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1703:139
  wire [31:0] _MUX1556__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1702:169
  wire        _GT1555__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1701:139
  wire [31:0] _dup1554__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1700:154
  wire [31:0] _dup1554__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1700:154
  wire [31:0] _dup1554__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1700:154
  wire [31:0] _SHR141553__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1699:97
  wire [31:0] _SUB1552__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1698:114
  wire [31:0] _MUX1550__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1696:169
  wire        _LT1549__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1695:139
  wire [31:0] _MUX1548__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1694:169
  wire        _GT1547__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1693:139
  wire [31:0] _dup1546__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1692:154
  wire [31:0] _dup1546__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1692:154
  wire [31:0] _dup1546__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1692:154
  wire [31:0] _SHR141545__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1691:97
  wire [31:0] _SUB1544__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1690:114
  wire [31:0] _MUX1542__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1688:169
  wire        _LT1541__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1687:139
  wire [31:0] _MUX1540__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1686:169
  wire        _GT1539__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1685:139
  wire [31:0] _dup1538__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1684:154
  wire [31:0] _dup1538__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1684:154
  wire [31:0] _dup1538__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1684:154
  wire [31:0] _SHR141537__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1683:97
  wire [31:0] _SUB1536__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1682:114
  wire [31:0] _MUX1534__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1680:169
  wire        _LT1533__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1679:139
  wire [31:0] _MUX1532__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1678:169
  wire        _GT1531__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1677:139
  wire [31:0] _dup1530__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1676:154
  wire [31:0] _dup1530__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1676:154
  wire [31:0] _dup1530__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1676:154
  wire [31:0] _SHR141529__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1675:97
  wire [31:0] _SUB1528__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1674:114
  wire [31:0] _MUX1526__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1672:169
  wire        _LT1525__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1671:139
  wire [31:0] _MUX1524__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1670:169
  wire        _GT1523__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1669:139
  wire [31:0] _dup1522__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1668:154
  wire [31:0] _dup1522__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1668:154
  wire [31:0] _dup1522__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1668:154
  wire [31:0] _SHR141521__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1667:97
  wire [31:0] _ADD1520__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1666:135
  wire [31:0] _dup1519__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1665:116
  wire [31:0] _dup1519__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1665:116
  wire [31:0] _dup1518__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1664:116
  wire [31:0] _dup1518__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1664:116
  wire [31:0] _MUX1516__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1662:169
  wire        _LT1515__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1661:139
  wire [31:0] _MUX1514__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1660:169
  wire        _GT1513__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1659:139
  wire [31:0] _dup1512__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1658:154
  wire [31:0] _dup1512__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1658:154
  wire [31:0] _dup1512__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1658:154
  wire [31:0] _SHR141511__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1657:97
  wire [31:0] _ADD1510__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1656:135
  wire [31:0] _dup1509__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1655:116
  wire [31:0] _dup1509__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1655:116
  wire [31:0] _dup1508__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1654:116
  wire [31:0] _dup1508__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1654:116
  wire [31:0] _MUX1506__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1652:169
  wire        _LT1505__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1651:139
  wire [31:0] _MUX1504__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1650:169
  wire        _GT1503__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1649:139
  wire [31:0] _dup1502__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1648:154
  wire [31:0] _dup1502__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1648:154
  wire [31:0] _dup1502__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1648:154
  wire [31:0] _SHR141501__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1647:97
  wire [31:0] _ADD1500__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1646:135
  wire [31:0] _dup1499__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1645:116
  wire [31:0] _dup1499__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1645:116
  wire [31:0] _dup1498__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1644:116
  wire [31:0] _dup1498__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1644:116
  wire [31:0] _MUX1496__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1642:169
  wire        _LT1495__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1641:139
  wire [31:0] _MUX1494__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1640:169
  wire        _GT1493__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1639:139
  wire [31:0] _dup1492__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1638:154
  wire [31:0] _dup1492__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1638:154
  wire [31:0] _dup1492__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1638:154
  wire [31:0] _SHR141491__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1637:97
  wire [31:0] _ADD1490__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1636:135
  wire [31:0] _dup1489__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1635:116
  wire [31:0] _dup1489__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1635:116
  wire [31:0] _dup1488__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1634:116
  wire [31:0] _dup1488__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1634:116
  wire [31:0] _SHR81487__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1633:91
  wire [31:0] _ADD1486__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1632:135
  wire [31:0] _MUL1485__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1631:136
  wire [31:0] _SUB1484__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1630:114
  wire [31:0] _SHR81483__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1629:91
  wire [31:0] _ADD1482__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1628:135
  wire [31:0] _MUL1481__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1627:136
  wire [31:0] _ADD1480__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1626:135
  wire [31:0] _dup1479__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1625:116
  wire [31:0] _dup1479__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1625:116
  wire [31:0] _dup1478__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1624:116
  wire [31:0] _dup1478__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1624:116
  wire [31:0] _SUB1477__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1623:114
  wire [31:0] _ADD1476__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1622:135
  wire [31:0] _dup1475__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1621:116
  wire [31:0] _dup1475__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1621:116
  wire [31:0] _dup1474__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1620:116
  wire [31:0] _dup1474__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1620:116
  wire [31:0] _SUB1473__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1619:114
  wire [31:0] _ADD1472__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1618:135
  wire [31:0] _dup1471__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1617:116
  wire [31:0] _dup1471__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1617:116
  wire [31:0] _dup1470__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1616:116
  wire [31:0] _dup1470__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1616:116
  wire [31:0] _SUB1469__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1615:114
  wire [31:0] _ADD1468__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1614:135
  wire [31:0] _dup1467__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1613:116
  wire [31:0] _dup1467__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1613:116
  wire [31:0] _dup1466__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1612:116
  wire [31:0] _dup1466__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1612:116
  wire [31:0] _SUB1465__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1611:114
  wire [31:0] _ADD1464__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1610:135
  wire [31:0] _dup1463__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1609:116
  wire [31:0] _dup1463__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1609:116
  wire [31:0] _dup1462__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1608:116
  wire [31:0] _dup1462__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1608:116
  wire [31:0] _SHR31461__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1607:93
  wire [31:0] _ADD1460__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1606:135
  wire [31:0] _MUL1459__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1605:136
  wire [31:0] _SHR31458__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1604:93
  wire [31:0] _SUB1457__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1603:114
  wire [31:0] _dup1456__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1602:116
  wire [31:0] _dup1456__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1602:116
  wire [31:0] _MUL1455__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1601:136
  wire [31:0] _ADD1454__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1600:135
  wire [31:0] _MUL1453__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1599:136
  wire [31:0] _ADD1452__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1598:135
  wire [31:0] _dup1451__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1597:116
  wire [31:0] _dup1451__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1597:116
  wire [31:0] _dup1450__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1596:116
  wire [31:0] _dup1450__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1596:116
  wire [31:0] _SUB1449__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1595:114
  wire [31:0] _ADD1448__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1594:135
  wire [31:0] _dup1447__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1593:116
  wire [31:0] _dup1447__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1593:116
  wire [31:0] _dup1446__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1592:116
  wire [31:0] _dup1446__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1592:116
  wire [31:0] _SHR31445__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1591:93
  wire [31:0] _SUB1444__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1590:114
  wire [31:0] _MUL1443__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1589:136
  wire [31:0] _SHR31442__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1588:93
  wire [31:0] _SUB1441__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1587:114
  wire [31:0] _dup1440__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1586:116
  wire [31:0] _dup1440__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1586:116
  wire [31:0] _MUL1439__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1585:136
  wire [31:0] _ADD1438__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1584:135
  wire [31:0] _MUL1437__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1583:136
  wire [31:0] _ADD1436__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1582:135
  wire [31:0] _dup1435__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1581:116
  wire [31:0] _dup1435__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1581:116
  wire [31:0] _dup1434__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1580:116
  wire [31:0] _dup1434__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1580:116
  wire [31:0] _SHR31433__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1579:93
  wire [31:0] _SUB1432__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1578:114
  wire [31:0] _MUL1431__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1577:136
  wire [31:0] _SHR31430__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1576:93
  wire [31:0] _ADD1429__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1575:135
  wire [31:0] _dup1428__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1574:116
  wire [31:0] _dup1428__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1574:116
  wire [31:0] _MUL1427__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1573:136
  wire [31:0] _ADD1426__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1572:135
  wire [31:0] _MUL1425__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1571:136
  wire [31:0] _ADD1424__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1570:135
  wire [31:0] _dup1423__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1569:116
  wire [31:0] _dup1423__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1569:116
  wire [31:0] _dup1422__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1568:116
  wire [31:0] _dup1422__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1568:116
  wire [31:0] _ADD1421__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1567:135
  wire [31:0] _SHL81420__dfc_wire_1923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1566:93
  wire [31:0] _CAST1419__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1565:88
  wire [31:0] _CAST1418__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1564:88
  wire [31:0] _CAST1417__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1563:88
  wire [31:0] _CAST1416__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1562:88
  wire [31:0] _CAST1415__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1561:88
  wire [31:0] _CAST1414__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1560:88
  wire [31:0] _CAST1413__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1559:88
  wire [31:0] _SHL81412__dfc_wire_1923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1558:93
  wire [31:0] _CAST1411__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1557:88
  wire [31:0] _MUX1409__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1555:169
  wire        _LT1408__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1554:139
  wire [31:0] _MUX1407__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1553:169
  wire        _GT1406__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1552:139
  wire [31:0] _dup1405__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1551:154
  wire [31:0] _dup1405__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1551:154
  wire [31:0] _dup1405__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1551:154
  wire [31:0] _SHR141404__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1550:97
  wire [31:0] _SUB1403__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1549:114
  wire [31:0] _MUX1401__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1547:169
  wire        _LT1400__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1546:139
  wire [31:0] _MUX1399__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1545:169
  wire        _GT1398__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1544:139
  wire [31:0] _dup1397__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1543:154
  wire [31:0] _dup1397__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1543:154
  wire [31:0] _dup1397__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1543:154
  wire [31:0] _SHR141396__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1542:97
  wire [31:0] _SUB1395__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1541:114
  wire [31:0] _MUX1393__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1539:169
  wire        _LT1392__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1538:139
  wire [31:0] _MUX1391__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1537:169
  wire        _GT1390__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1536:139
  wire [31:0] _dup1389__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1535:154
  wire [31:0] _dup1389__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1535:154
  wire [31:0] _dup1389__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1535:154
  wire [31:0] _SHR141388__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1534:97
  wire [31:0] _SUB1387__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1533:114
  wire [31:0] _MUX1385__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1531:169
  wire        _LT1384__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1530:139
  wire [31:0] _MUX1383__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1529:169
  wire        _GT1382__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1528:139
  wire [31:0] _dup1381__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1527:154
  wire [31:0] _dup1381__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1527:154
  wire [31:0] _dup1381__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1527:154
  wire [31:0] _SHR141380__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1526:97
  wire [31:0] _SUB1379__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1525:114
  wire [31:0] _MUX1377__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1523:169
  wire        _LT1376__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1522:139
  wire [31:0] _MUX1375__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1521:169
  wire        _GT1374__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1520:139
  wire [31:0] _dup1373__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1519:154
  wire [31:0] _dup1373__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1519:154
  wire [31:0] _dup1373__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1519:154
  wire [31:0] _SHR141372__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1518:97
  wire [31:0] _ADD1371__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1517:135
  wire [31:0] _dup1370__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1516:116
  wire [31:0] _dup1370__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1516:116
  wire [31:0] _dup1369__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1515:116
  wire [31:0] _dup1369__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1515:116
  wire [31:0] _MUX1367__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1513:169
  wire        _LT1366__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1512:139
  wire [31:0] _MUX1365__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1511:169
  wire        _GT1364__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1510:139
  wire [31:0] _dup1363__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1509:154
  wire [31:0] _dup1363__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1509:154
  wire [31:0] _dup1363__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1509:154
  wire [31:0] _SHR141362__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1508:97
  wire [31:0] _ADD1361__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1507:135
  wire [31:0] _dup1360__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1506:116
  wire [31:0] _dup1360__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1506:116
  wire [31:0] _dup1359__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1505:116
  wire [31:0] _dup1359__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1505:116
  wire [31:0] _MUX1357__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1503:169
  wire        _LT1356__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1502:139
  wire [31:0] _MUX1355__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1501:169
  wire        _GT1354__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1500:139
  wire [31:0] _dup1353__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1499:154
  wire [31:0] _dup1353__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1499:154
  wire [31:0] _dup1353__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1499:154
  wire [31:0] _SHR141352__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1498:97
  wire [31:0] _ADD1351__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1497:135
  wire [31:0] _dup1350__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1496:116
  wire [31:0] _dup1350__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1496:116
  wire [31:0] _dup1349__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1495:116
  wire [31:0] _dup1349__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1495:116
  wire [31:0] _MUX1347__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1493:169
  wire        _LT1346__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1492:139
  wire [31:0] _MUX1345__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1491:169
  wire        _GT1344__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1490:139
  wire [31:0] _dup1343__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1489:154
  wire [31:0] _dup1343__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1489:154
  wire [31:0] _dup1343__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1489:154
  wire [31:0] _SHR141342__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1488:97
  wire [31:0] _ADD1341__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1487:135
  wire [31:0] _dup1340__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1486:116
  wire [31:0] _dup1340__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1486:116
  wire [31:0] _dup1339__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1485:116
  wire [31:0] _dup1339__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1485:116
  wire [31:0] _SHR81338__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1484:91
  wire [31:0] _ADD1337__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1483:135
  wire [31:0] _MUL1336__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1482:136
  wire [31:0] _SUB1335__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1481:114
  wire [31:0] _SHR81334__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1480:91
  wire [31:0] _ADD1333__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1479:135
  wire [31:0] _MUL1332__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1478:136
  wire [31:0] _ADD1331__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1477:135
  wire [31:0] _dup1330__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1476:116
  wire [31:0] _dup1330__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1476:116
  wire [31:0] _dup1329__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1475:116
  wire [31:0] _dup1329__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1475:116
  wire [31:0] _SUB1328__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1474:114
  wire [31:0] _ADD1327__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1473:135
  wire [31:0] _dup1326__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1472:116
  wire [31:0] _dup1326__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1472:116
  wire [31:0] _dup1325__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1471:116
  wire [31:0] _dup1325__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1471:116
  wire [31:0] _SUB1324__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1470:114
  wire [31:0] _ADD1323__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1469:135
  wire [31:0] _dup1322__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1468:116
  wire [31:0] _dup1322__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1468:116
  wire [31:0] _dup1321__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1467:116
  wire [31:0] _dup1321__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1467:116
  wire [31:0] _SUB1320__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1466:114
  wire [31:0] _ADD1319__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1465:135
  wire [31:0] _dup1318__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1464:116
  wire [31:0] _dup1318__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1464:116
  wire [31:0] _dup1317__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1463:116
  wire [31:0] _dup1317__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1463:116
  wire [31:0] _SUB1316__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1462:114
  wire [31:0] _ADD1315__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1461:135
  wire [31:0] _dup1314__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1460:116
  wire [31:0] _dup1314__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1460:116
  wire [31:0] _dup1313__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1459:116
  wire [31:0] _dup1313__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1459:116
  wire [31:0] _SHR31312__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1458:93
  wire [31:0] _ADD1311__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1457:135
  wire [31:0] _MUL1310__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1456:136
  wire [31:0] _SHR31309__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1455:93
  wire [31:0] _SUB1308__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1454:114
  wire [31:0] _dup1307__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1453:116
  wire [31:0] _dup1307__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1453:116
  wire [31:0] _MUL1306__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1452:136
  wire [31:0] _ADD1305__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1451:135
  wire [31:0] _MUL1304__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1450:136
  wire [31:0] _ADD1303__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1449:135
  wire [31:0] _dup1302__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1448:116
  wire [31:0] _dup1302__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1448:116
  wire [31:0] _dup1301__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1447:116
  wire [31:0] _dup1301__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1447:116
  wire [31:0] _SUB1300__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1446:114
  wire [31:0] _ADD1299__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1445:135
  wire [31:0] _dup1298__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1444:116
  wire [31:0] _dup1298__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1444:116
  wire [31:0] _dup1297__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1443:116
  wire [31:0] _dup1297__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1443:116
  wire [31:0] _SHR31296__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1442:93
  wire [31:0] _SUB1295__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1441:114
  wire [31:0] _MUL1294__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1440:136
  wire [31:0] _SHR31293__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1439:93
  wire [31:0] _SUB1292__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1438:114
  wire [31:0] _dup1291__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1437:116
  wire [31:0] _dup1291__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1437:116
  wire [31:0] _MUL1290__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1436:136
  wire [31:0] _ADD1289__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1435:135
  wire [31:0] _MUL1288__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1434:136
  wire [31:0] _ADD1287__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1433:135
  wire [31:0] _dup1286__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1432:116
  wire [31:0] _dup1286__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1432:116
  wire [31:0] _dup1285__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1431:116
  wire [31:0] _dup1285__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1431:116
  wire [31:0] _SHR31284__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1430:93
  wire [31:0] _SUB1283__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1429:114
  wire [31:0] _MUL1282__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1428:136
  wire [31:0] _SHR31281__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1427:93
  wire [31:0] _ADD1280__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1426:135
  wire [31:0] _dup1279__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1425:116
  wire [31:0] _dup1279__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1425:116
  wire [31:0] _MUL1278__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1424:136
  wire [31:0] _ADD1277__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1423:135
  wire [31:0] _MUL1276__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1422:136
  wire [31:0] _ADD1275__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1421:135
  wire [31:0] _dup1274__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1420:116
  wire [31:0] _dup1274__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1420:116
  wire [31:0] _dup1273__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1419:116
  wire [31:0] _dup1273__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1419:116
  wire [31:0] _ADD1272__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1418:135
  wire [31:0] _SHL81271__dfc_wire_1923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1417:93
  wire [31:0] _CAST1270__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1416:88
  wire [31:0] _CAST1269__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1415:88
  wire [31:0] _CAST1268__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1414:88
  wire [31:0] _CAST1267__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1413:88
  wire [31:0] _CAST1266__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1412:88
  wire [31:0] _CAST1265__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1411:88
  wire [31:0] _CAST1264__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1410:88
  wire [31:0] _SHL81263__dfc_wire_1923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1409:93
  wire [31:0] _CAST1262__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1408:88
  wire [31:0] _MUX1260__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1406:169
  wire        _LT1259__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1405:139
  wire [31:0] _MUX1258__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1404:169
  wire        _GT1257__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1403:139
  wire [31:0] _dup1256__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1402:154
  wire [31:0] _dup1256__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1402:154
  wire [31:0] _dup1256__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1402:154
  wire [31:0] _SHR141255__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1401:97
  wire [31:0] _SUB1254__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1400:114
  wire [31:0] _MUX1252__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1398:169
  wire        _LT1251__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1397:139
  wire [31:0] _MUX1250__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1396:169
  wire        _GT1249__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1395:139
  wire [31:0] _dup1248__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1394:154
  wire [31:0] _dup1248__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1394:154
  wire [31:0] _dup1248__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1394:154
  wire [31:0] _SHR141247__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1393:97
  wire [31:0] _SUB1246__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1392:114
  wire [31:0] _MUX1244__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1390:169
  wire        _LT1243__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1389:139
  wire [31:0] _MUX1242__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1388:169
  wire        _GT1241__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1387:139
  wire [31:0] _dup1240__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1386:154
  wire [31:0] _dup1240__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1386:154
  wire [31:0] _dup1240__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1386:154
  wire [31:0] _SHR141239__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1385:97
  wire [31:0] _SUB1238__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1384:114
  wire [31:0] _MUX1236__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1382:169
  wire        _LT1235__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1381:139
  wire [31:0] _MUX1234__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1380:169
  wire        _GT1233__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1379:139
  wire [31:0] _dup1232__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1378:154
  wire [31:0] _dup1232__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1378:154
  wire [31:0] _dup1232__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1378:154
  wire [31:0] _SHR141231__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1377:97
  wire [31:0] _SUB1230__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1376:114
  wire [31:0] _MUX1228__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1374:169
  wire        _LT1227__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1373:139
  wire [31:0] _MUX1226__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1372:169
  wire        _GT1225__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1371:139
  wire [31:0] _dup1224__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1370:154
  wire [31:0] _dup1224__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1370:154
  wire [31:0] _dup1224__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1370:154
  wire [31:0] _SHR141223__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1369:97
  wire [31:0] _ADD1222__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1368:135
  wire [31:0] _dup1221__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1367:116
  wire [31:0] _dup1221__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1367:116
  wire [31:0] _dup1220__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1366:116
  wire [31:0] _dup1220__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1366:116
  wire [31:0] _MUX1218__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1364:169
  wire        _LT1217__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1363:139
  wire [31:0] _MUX1216__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1362:169
  wire        _GT1215__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1361:139
  wire [31:0] _dup1214__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1360:154
  wire [31:0] _dup1214__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1360:154
  wire [31:0] _dup1214__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1360:154
  wire [31:0] _SHR141213__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1359:97
  wire [31:0] _ADD1212__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1358:135
  wire [31:0] _dup1211__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1357:116
  wire [31:0] _dup1211__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1357:116
  wire [31:0] _dup1210__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1356:116
  wire [31:0] _dup1210__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1356:116
  wire [31:0] _MUX1208__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1354:169
  wire        _LT1207__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1353:139
  wire [31:0] _MUX1206__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1352:169
  wire        _GT1205__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1351:139
  wire [31:0] _dup1204__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1350:154
  wire [31:0] _dup1204__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1350:154
  wire [31:0] _dup1204__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1350:154
  wire [31:0] _SHR141203__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1349:97
  wire [31:0] _ADD1202__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1348:135
  wire [31:0] _dup1201__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1347:116
  wire [31:0] _dup1201__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1347:116
  wire [31:0] _dup1200__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1346:116
  wire [31:0] _dup1200__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1346:116
  wire [31:0] _MUX1198__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1344:169
  wire        _LT1197__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1343:139
  wire [31:0] _MUX1196__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1342:169
  wire        _GT1195__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1341:139
  wire [31:0] _dup1194__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1340:154
  wire [31:0] _dup1194__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1340:154
  wire [31:0] _dup1194__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1340:154
  wire [31:0] _SHR141193__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1339:97
  wire [31:0] _ADD1192__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1338:135
  wire [31:0] _dup1191__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1337:116
  wire [31:0] _dup1191__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1337:116
  wire [31:0] _dup1190__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1336:116
  wire [31:0] _dup1190__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1336:116
  wire [31:0] _SHR81189__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1335:91
  wire [31:0] _ADD1188__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1334:135
  wire [31:0] _MUL1187__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1333:136
  wire [31:0] _SUB1186__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1332:114
  wire [31:0] _SHR81185__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1331:91
  wire [31:0] _ADD1184__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1330:135
  wire [31:0] _MUL1183__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1329:136
  wire [31:0] _ADD1182__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1328:135
  wire [31:0] _dup1181__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1327:116
  wire [31:0] _dup1181__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1327:116
  wire [31:0] _dup1180__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1326:116
  wire [31:0] _dup1180__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1326:116
  wire [31:0] _SUB1179__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1325:114
  wire [31:0] _ADD1178__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1324:135
  wire [31:0] _dup1177__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1323:116
  wire [31:0] _dup1177__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1323:116
  wire [31:0] _dup1176__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1322:116
  wire [31:0] _dup1176__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1322:116
  wire [31:0] _SUB1175__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1321:114
  wire [31:0] _ADD1174__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1320:135
  wire [31:0] _dup1173__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1319:116
  wire [31:0] _dup1173__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1319:116
  wire [31:0] _dup1172__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1318:116
  wire [31:0] _dup1172__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1318:116
  wire [31:0] _SUB1171__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1317:114
  wire [31:0] _ADD1170__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1316:135
  wire [31:0] _dup1169__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1315:116
  wire [31:0] _dup1169__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1315:116
  wire [31:0] _dup1168__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1314:116
  wire [31:0] _dup1168__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1314:116
  wire [31:0] _SUB1167__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1313:114
  wire [31:0] _ADD1166__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1312:135
  wire [31:0] _dup1165__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1311:116
  wire [31:0] _dup1165__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1311:116
  wire [31:0] _dup1164__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1310:116
  wire [31:0] _dup1164__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1310:116
  wire [31:0] _SHR31163__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1309:93
  wire [31:0] _ADD1162__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1308:135
  wire [31:0] _MUL1161__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1307:136
  wire [31:0] _SHR31160__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1306:93
  wire [31:0] _SUB1159__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1305:114
  wire [31:0] _dup1158__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1304:116
  wire [31:0] _dup1158__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1304:116
  wire [31:0] _MUL1157__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1303:136
  wire [31:0] _ADD1156__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1302:135
  wire [31:0] _MUL1155__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1301:136
  wire [31:0] _ADD1154__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1300:135
  wire [31:0] _dup1153__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1299:116
  wire [31:0] _dup1153__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1299:116
  wire [31:0] _dup1152__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1298:116
  wire [31:0] _dup1152__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1298:116
  wire [31:0] _SUB1151__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1297:114
  wire [31:0] _ADD1150__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1296:135
  wire [31:0] _dup1149__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1295:116
  wire [31:0] _dup1149__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1295:116
  wire [31:0] _dup1148__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1294:116
  wire [31:0] _dup1148__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1294:116
  wire [31:0] _SHR31147__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1293:93
  wire [31:0] _SUB1146__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1292:114
  wire [31:0] _MUL1145__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1291:136
  wire [31:0] _SHR31144__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1290:93
  wire [31:0] _SUB1143__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1289:114
  wire [31:0] _dup1142__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1288:116
  wire [31:0] _dup1142__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1288:116
  wire [31:0] _MUL1141__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1287:136
  wire [31:0] _ADD1140__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1286:135
  wire [31:0] _MUL1139__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1285:136
  wire [31:0] _ADD1138__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1284:135
  wire [31:0] _dup1137__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1283:116
  wire [31:0] _dup1137__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1283:116
  wire [31:0] _dup1136__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1282:116
  wire [31:0] _dup1136__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1282:116
  wire [31:0] _SHR31135__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1281:93
  wire [31:0] _SUB1134__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1280:114
  wire [31:0] _MUL1133__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1279:136
  wire [31:0] _SHR31132__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1278:93
  wire [31:0] _ADD1131__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1277:135
  wire [31:0] _dup1130__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1276:116
  wire [31:0] _dup1130__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1276:116
  wire [31:0] _MUL1129__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1275:136
  wire [31:0] _ADD1128__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1274:135
  wire [31:0] _MUL1127__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1273:136
  wire [31:0] _ADD1126__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1272:135
  wire [31:0] _dup1125__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1271:116
  wire [31:0] _dup1125__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1271:116
  wire [31:0] _dup1124__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1270:116
  wire [31:0] _dup1124__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1270:116
  wire [31:0] _ADD1123__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1269:135
  wire [31:0] _SHL81122__dfc_wire_1923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1268:93
  wire [31:0] _CAST1121__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1267:88
  wire [31:0] _CAST1120__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1266:88
  wire [31:0] _CAST1119__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1265:88
  wire [31:0] _CAST1118__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1264:88
  wire [31:0] _CAST1117__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1263:88
  wire [31:0] _CAST1116__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1262:88
  wire [31:0] _CAST1115__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1261:88
  wire [31:0] _SHL81114__dfc_wire_1923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1260:93
  wire [31:0] _CAST1113__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1259:88
  wire [31:0] _MUX1111__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1257:169
  wire        _LT1110__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1256:139
  wire [31:0] _MUX1109__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1255:169
  wire        _GT1108__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1254:139
  wire [31:0] _dup1107__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1253:154
  wire [31:0] _dup1107__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1253:154
  wire [31:0] _dup1107__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1253:154
  wire [31:0] _SHR141106__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1252:97
  wire [31:0] _SUB1105__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1251:114
  wire [31:0] _MUX1103__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1249:169
  wire        _LT1102__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1248:139
  wire [31:0] _MUX1101__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1247:169
  wire        _GT1100__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1246:139
  wire [31:0] _dup1099__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1245:154
  wire [31:0] _dup1099__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1245:154
  wire [31:0] _dup1099__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1245:154
  wire [31:0] _SHR141098__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1244:97
  wire [31:0] _SUB1097__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1243:114
  wire [31:0] _MUX1095__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1241:169
  wire        _LT1094__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1240:139
  wire [31:0] _MUX1093__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1239:169
  wire        _GT1092__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1238:139
  wire [31:0] _dup1091__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1237:154
  wire [31:0] _dup1091__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1237:154
  wire [31:0] _dup1091__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1237:154
  wire [31:0] _SHR141090__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1236:97
  wire [31:0] _SUB1089__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1235:114
  wire [31:0] _MUX1087__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1233:169
  wire        _LT1086__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1232:139
  wire [31:0] _MUX1085__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1231:169
  wire        _GT1084__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1230:139
  wire [31:0] _dup1083__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1229:154
  wire [31:0] _dup1083__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1229:154
  wire [31:0] _dup1083__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1229:154
  wire [31:0] _SHR141082__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1228:97
  wire [31:0] _SUB1081__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1227:114
  wire [31:0] _MUX1079__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1225:169
  wire        _LT1078__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1224:139
  wire [31:0] _MUX1077__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1223:169
  wire        _GT1076__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1222:139
  wire [31:0] _dup1075__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1221:154
  wire [31:0] _dup1075__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1221:154
  wire [31:0] _dup1075__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1221:154
  wire [31:0] _SHR141074__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1220:97
  wire [31:0] _ADD1073__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1219:135
  wire [31:0] _dup1072__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1218:116
  wire [31:0] _dup1072__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1218:116
  wire [31:0] _dup1071__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1217:116
  wire [31:0] _dup1071__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1217:116
  wire [31:0] _MUX1069__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1215:169
  wire        _LT1068__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1214:139
  wire [31:0] _MUX1067__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1213:169
  wire        _GT1066__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1212:139
  wire [31:0] _dup1065__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1211:154
  wire [31:0] _dup1065__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1211:154
  wire [31:0] _dup1065__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1211:154
  wire [31:0] _SHR141064__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1210:97
  wire [31:0] _ADD1063__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1209:135
  wire [31:0] _dup1062__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1208:116
  wire [31:0] _dup1062__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1208:116
  wire [31:0] _dup1061__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1207:116
  wire [31:0] _dup1061__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1207:116
  wire [31:0] _MUX1059__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1205:169
  wire        _LT1058__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1204:139
  wire [31:0] _MUX1057__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1203:169
  wire        _GT1056__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1202:139
  wire [31:0] _dup1055__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1201:154
  wire [31:0] _dup1055__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1201:154
  wire [31:0] _dup1055__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1201:154
  wire [31:0] _SHR141054__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1200:97
  wire [31:0] _ADD1053__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1199:135
  wire [31:0] _dup1052__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1198:116
  wire [31:0] _dup1052__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1198:116
  wire [31:0] _dup1051__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1197:116
  wire [31:0] _dup1051__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1197:116
  wire [31:0] _MUX1049__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1195:169
  wire        _LT1048__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1194:139
  wire [31:0] _MUX1047__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1193:169
  wire        _GT1046__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1192:139
  wire [31:0] _dup1045__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1191:154
  wire [31:0] _dup1045__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1191:154
  wire [31:0] _dup1045__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1191:154
  wire [31:0] _SHR141044__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1190:97
  wire [31:0] _ADD1043__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1189:135
  wire [31:0] _dup1042__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1188:116
  wire [31:0] _dup1042__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1188:116
  wire [31:0] _dup1041__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1187:116
  wire [31:0] _dup1041__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1187:116
  wire [31:0] _SHR81040__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1186:91
  wire [31:0] _ADD1039__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1185:135
  wire [31:0] _MUL1038__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1184:136
  wire [31:0] _SUB1037__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1183:114
  wire [31:0] _SHR81036__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1182:91
  wire [31:0] _ADD1035__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1181:135
  wire [31:0] _MUL1034__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1180:136
  wire [31:0] _ADD1033__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1179:135
  wire [31:0] _dup1032__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1178:116
  wire [31:0] _dup1032__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1178:116
  wire [31:0] _dup1031__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1177:116
  wire [31:0] _dup1031__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1177:116
  wire [31:0] _SUB1030__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1176:114
  wire [31:0] _ADD1029__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1175:135
  wire [31:0] _dup1028__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1174:116
  wire [31:0] _dup1028__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1174:116
  wire [31:0] _dup1027__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1173:116
  wire [31:0] _dup1027__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1173:116
  wire [31:0] _SUB1026__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1172:114
  wire [31:0] _ADD1025__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1171:135
  wire [31:0] _dup1024__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1170:116
  wire [31:0] _dup1024__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1170:116
  wire [31:0] _dup1023__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1169:116
  wire [31:0] _dup1023__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1169:116
  wire [31:0] _SUB1022__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1168:114
  wire [31:0] _ADD1021__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1167:135
  wire [31:0] _dup1020__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1166:116
  wire [31:0] _dup1020__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1166:116
  wire [31:0] _dup1019__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1165:116
  wire [31:0] _dup1019__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1165:116
  wire [31:0] _SUB1018__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1164:114
  wire [31:0] _ADD1017__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1163:135
  wire [31:0] _dup1016__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1162:116
  wire [31:0] _dup1016__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1162:116
  wire [31:0] _dup1015__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1161:116
  wire [31:0] _dup1015__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1161:116
  wire [31:0] _SHR31014__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1160:93
  wire [31:0] _ADD1013__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1159:135
  wire [31:0] _MUL1012__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1158:136
  wire [31:0] _SHR31011__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1157:93
  wire [31:0] _SUB1010__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1156:114
  wire [31:0] _dup1009__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1155:116
  wire [31:0] _dup1009__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1155:116
  wire [31:0] _MUL1008__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1154:136
  wire [31:0] _ADD1007__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1153:135
  wire [31:0] _MUL1006__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1152:136
  wire [31:0] _ADD1005__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1151:135
  wire [31:0] _dup1004__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1150:116
  wire [31:0] _dup1004__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1150:116
  wire [31:0] _dup1003__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1149:116
  wire [31:0] _dup1003__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1149:116
  wire [31:0] _SUB1002__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1148:114
  wire [31:0] _ADD1001__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1147:135
  wire [31:0] _dup1000__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1146:116
  wire [31:0] _dup1000__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1146:116
  wire [31:0] _dup999__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1145:111
  wire [31:0] _dup999__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1145:111
  wire [31:0] _SHR3998__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1144:89
  wire [31:0] _SUB997__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1143:109
  wire [31:0] _MUL996__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1142:131
  wire [31:0] _SHR3995__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1141:89
  wire [31:0] _SUB994__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1140:109
  wire [31:0] _dup993__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1139:111
  wire [31:0] _dup993__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1139:111
  wire [31:0] _MUL992__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1138:131
  wire [31:0] _ADD991__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1137:130
  wire [31:0] _MUL990__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1136:131
  wire [31:0] _ADD989__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1135:130
  wire [31:0] _dup988__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1134:111
  wire [31:0] _dup988__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1134:111
  wire [31:0] _dup987__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1133:111
  wire [31:0] _dup987__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1133:111
  wire [31:0] _SHR3986__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1132:89
  wire [31:0] _SUB985__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1131:109
  wire [31:0] _MUL984__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1130:131
  wire [31:0] _SHR3983__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1129:89
  wire [31:0] _ADD982__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1128:130
  wire [31:0] _dup981__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1127:111
  wire [31:0] _dup981__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1127:111
  wire [31:0] _MUL980__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1126:131
  wire [31:0] _ADD979__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1125:130
  wire [31:0] _MUL978__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1124:131
  wire [31:0] _ADD977__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1123:130
  wire [31:0] _dup976__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1122:111
  wire [31:0] _dup976__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1122:111
  wire [31:0] _dup975__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1121:111
  wire [31:0] _dup975__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1121:111
  wire [31:0] _ADD974__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1120:130
  wire [31:0] _SHL8973__dfc_wire_1923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1119:89
  wire [31:0] _CAST972__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1118:84
  wire [31:0] _CAST971__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1117:84
  wire [31:0] _CAST970__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1116:84
  wire [31:0] _CAST969__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1115:84
  wire [31:0] _CAST968__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1114:84
  wire [31:0] _CAST967__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1113:84
  wire [31:0] _CAST966__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1112:84
  wire [31:0] _SHL8965__dfc_wire_1923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1111:89
  wire [31:0] _CAST964__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1110:84
  wire [31:0] _MUX962__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1108:163
  wire        _LT961__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1107:134
  wire [31:0] _MUX960__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1106:163
  wire        _GT959__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1105:134
  wire [31:0] _dup958__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1104:148
  wire [31:0] _dup958__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1104:148
  wire [31:0] _dup958__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1104:148
  wire [31:0] _SHR14957__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1103:93
  wire [31:0] _SUB956__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1102:109
  wire [31:0] _MUX954__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1100:163
  wire        _LT953__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1099:134
  wire [31:0] _MUX952__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1098:163
  wire        _GT951__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1097:134
  wire [31:0] _dup950__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1096:148
  wire [31:0] _dup950__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1096:148
  wire [31:0] _dup950__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1096:148
  wire [31:0] _SHR14949__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1095:93
  wire [31:0] _SUB948__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1094:109
  wire [31:0] _MUX946__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1092:163
  wire        _LT945__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1091:134
  wire [31:0] _MUX944__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1090:163
  wire        _GT943__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1089:134
  wire [31:0] _dup942__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1088:148
  wire [31:0] _dup942__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1088:148
  wire [31:0] _dup942__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1088:148
  wire [31:0] _SHR14941__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1087:93
  wire [31:0] _SUB940__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1086:109
  wire [31:0] _MUX938__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1084:163
  wire        _LT937__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1083:134
  wire [31:0] _MUX936__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1082:163
  wire        _GT935__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1081:134
  wire [31:0] _dup934__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1080:148
  wire [31:0] _dup934__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1080:148
  wire [31:0] _dup934__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1080:148
  wire [31:0] _SHR14933__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1079:93
  wire [31:0] _SUB932__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1078:109
  wire [31:0] _MUX930__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1076:163
  wire        _LT929__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1075:134
  wire [31:0] _MUX928__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1074:163
  wire        _GT927__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1073:134
  wire [31:0] _dup926__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1072:148
  wire [31:0] _dup926__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1072:148
  wire [31:0] _dup926__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1072:148
  wire [31:0] _SHR14925__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1071:93
  wire [31:0] _ADD924__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1070:130
  wire [31:0] _dup923__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1069:111
  wire [31:0] _dup923__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1069:111
  wire [31:0] _dup922__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1068:111
  wire [31:0] _dup922__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1068:111
  wire [31:0] _MUX920__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1066:163
  wire        _LT919__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1065:134
  wire [31:0] _MUX918__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1064:163
  wire        _GT917__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1063:134
  wire [31:0] _dup916__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1062:148
  wire [31:0] _dup916__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1062:148
  wire [31:0] _dup916__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1062:148
  wire [31:0] _SHR14915__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1061:93
  wire [31:0] _ADD914__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1060:130
  wire [31:0] _dup913__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1059:111
  wire [31:0] _dup913__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1059:111
  wire [31:0] _dup912__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1058:111
  wire [31:0] _dup912__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1058:111
  wire [31:0] _MUX910__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1056:163
  wire        _LT909__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1055:134
  wire [31:0] _MUX908__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1054:163
  wire        _GT907__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1053:134
  wire [31:0] _dup906__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1052:148
  wire [31:0] _dup906__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1052:148
  wire [31:0] _dup906__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1052:148
  wire [31:0] _SHR14905__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1051:93
  wire [31:0] _ADD904__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1050:130
  wire [31:0] _dup903__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1049:111
  wire [31:0] _dup903__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1049:111
  wire [31:0] _dup902__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1048:111
  wire [31:0] _dup902__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1048:111
  wire [31:0] _MUX900__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1046:163
  wire        _LT899__dfc_wire_2112;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1045:134
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2111;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2129;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2133;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2151;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2155;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2173;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2177;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2195;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2199;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2217;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2221;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2239;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2243;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2261;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2265;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2471;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2475;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2493;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2497;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2515;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2519;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2537;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2541;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2559;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2563;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2581;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2585;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2603;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2607;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2625;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2629;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2835;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2839;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2857;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2861;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2879;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2883;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2901;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2905;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2927;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2945;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2949;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2967;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2971;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2989;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_2993;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3199;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3203;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3221;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3225;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3243;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3247;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3265;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3269;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3287;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3291;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3309;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3313;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3331;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3335;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3353;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3357;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3563;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3567;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3585;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3589;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3607;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3611;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3629;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3633;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3651;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3655;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3673;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3677;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3695;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3699;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3717;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3721;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3927;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3931;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3949;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3953;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3971;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3975;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3993;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_3997;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4015;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4019;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4037;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4041;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4059;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4063;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4081;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4085;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4291;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4295;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4313;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4317;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4335;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4339;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4357;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4361;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4379;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4383;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4401;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4405;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4423;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4427;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4445;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4449;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4655;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4659;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4677;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4681;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4699;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4703;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4721;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4725;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4743;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4747;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4765;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4769;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4787;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4791;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4809;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _dup898_const_fix_32_0_1__00000000000000ff_4813;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
  wire [31:0] _MUX897__dfc_wire_2108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1043:163
  wire        _GT896__dfc_wire_2105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1042:134
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2111;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2129;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2133;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2151;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2155;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2173;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2177;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2195;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2199;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2217;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2221;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2239;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2243;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2261;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2265;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2471;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2475;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2493;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2497;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2515;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2519;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2537;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2541;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2559;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2563;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2581;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2585;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2603;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2607;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2625;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2629;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2835;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2839;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2857;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2861;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2879;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2883;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2901;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2905;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2927;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2945;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2949;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2967;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2971;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2989;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_2993;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3199;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3203;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3221;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3225;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3243;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3247;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3265;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3269;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3287;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3291;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3309;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3313;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3331;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3335;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3353;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3357;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3563;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3567;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3585;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3589;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3607;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3611;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3629;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3633;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3651;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3655;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3673;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3677;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3695;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3699;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3717;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3721;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3927;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3931;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3949;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3953;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3971;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3975;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3993;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_3997;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4015;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4019;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4037;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4041;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4059;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4063;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4081;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4085;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4291;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4295;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4313;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4317;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4335;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4339;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4357;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4361;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4379;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4383;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4401;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4405;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4423;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4427;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4445;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4449;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4655;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4659;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4677;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4681;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4699;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4703;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4721;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4725;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4743;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4747;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4765;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4769;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4787;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4791;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4809;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup895_const_fix_32_0_1__00000000000000ff_4813;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
  wire [31:0] _dup894__dfc_wire_2103_2106;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1040:148
  wire [31:0] _dup894__dfc_wire_2103_2110;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1040:148
  wire [31:0] _dup894__dfc_wire_2103_2113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1040:148
  wire [31:0] _SHR14893__dfc_wire_2103;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1039:93
  wire [31:0] _ADD892__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1038:130
  wire [31:0] _dup891__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1037:111
  wire [31:0] _dup891__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1037:111
  wire [31:0] _dup890__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1036:111
  wire [31:0] _dup890__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1036:111
  wire [31:0] _SHR8889__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1035:87
  wire [31:0] _ADD888__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1034:130
  wire [31:0] _MUL887__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1033:131
  wire [31:0] _SUB886__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1032:109
  wire [31:0] _SHR8885__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1031:87
  wire [31:0] _ADD884__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1030:130
  wire [31:0] _MUL883__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1029:131
  wire [31:0] _ADD882__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1028:130
  wire [31:0] _dup881__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1027:111
  wire [31:0] _dup881__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1027:111
  wire [31:0] _dup880__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1026:111
  wire [31:0] _dup880__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1026:111
  wire [31:0] _SUB879__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1025:109
  wire [31:0] _ADD878__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1024:130
  wire [31:0] _dup877__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1023:111
  wire [31:0] _dup877__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1023:111
  wire [31:0] _dup876__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1022:111
  wire [31:0] _dup876__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1022:111
  wire [31:0] _SUB875__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1021:109
  wire [31:0] _ADD874__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1020:130
  wire [31:0] _dup873__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1019:111
  wire [31:0] _dup873__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1019:111
  wire [31:0] _dup872__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1018:111
  wire [31:0] _dup872__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1018:111
  wire [31:0] _SUB871__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1017:109
  wire [31:0] _ADD870__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1016:130
  wire [31:0] _dup869__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1015:111
  wire [31:0] _dup869__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1015:111
  wire [31:0] _dup868__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1014:111
  wire [31:0] _dup868__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1014:111
  wire [31:0] _SUB867__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1013:109
  wire [31:0] _ADD866__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1012:130
  wire [31:0] _dup865__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1011:111
  wire [31:0] _dup865__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1011:111
  wire [31:0] _dup864__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1010:111
  wire [31:0] _dup864__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1010:111
  wire [31:0] _SHR3863__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1009:89
  wire [31:0] _ADD862__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1008:130
  wire [31:0] _MUL861__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1007:131
  wire [31:0] _SHR3860__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1006:89
  wire [31:0] _SUB859__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1005:109
  wire [31:0] _dup858__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1004:111
  wire [31:0] _dup858__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1004:111
  wire [31:0] _MUL857__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1003:131
  wire [31:0] _ADD856__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1002:130
  wire [31:0] _MUL855__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1001:131
  wire [31:0] _ADD854__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1000:130
  wire [31:0] _dup853__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:999:111
  wire [31:0] _dup853__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:999:111
  wire [31:0] _dup852__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:998:111
  wire [31:0] _dup852__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:998:111
  wire [31:0] _SUB851__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:997:109
  wire [31:0] _ADD850__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:996:130
  wire [31:0] _dup849__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:995:111
  wire [31:0] _dup849__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:995:111
  wire [31:0] _dup848__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:994:111
  wire [31:0] _dup848__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:994:111
  wire [31:0] _SHR3847__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:993:89
  wire [31:0] _SUB846__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:992:109
  wire [31:0] _MUL845__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:991:131
  wire [31:0] _SHR3844__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:990:89
  wire [31:0] _SUB843__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:989:109
  wire [31:0] _dup842__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:988:111
  wire [31:0] _dup842__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:988:111
  wire [31:0] _MUL841__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:987:131
  wire [31:0] _ADD840__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:986:130
  wire [31:0] _MUL839__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:985:131
  wire [31:0] _ADD838__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:984:130
  wire [31:0] _dup837__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:983:111
  wire [31:0] _dup837__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:983:111
  wire [31:0] _dup836__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:982:111
  wire [31:0] _dup836__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:982:111
  wire [31:0] _SHR3835__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:981:89
  wire [31:0] _SUB834__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:980:109
  wire [31:0] _MUL833__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:979:131
  wire [31:0] _SHR3832__dfc_wire_1968;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:978:89
  wire [31:0] _ADD831__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:977:130
  wire [31:0] _dup830__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:976:111
  wire [31:0] _dup830__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:976:111
  wire [31:0] _MUL829__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:975:131
  wire [31:0] _ADD828__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:974:130
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_1960;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_1988;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_2024;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_2324;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_2352;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_2388;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_2688;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_2716;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_2752;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_3052;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_3080;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_3116;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_3416;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_3444;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_3480;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_3780;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_3808;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_3844;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_4144;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_4172;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_4208;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_4508;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_4536;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _dup827_const_fix_32_0_1__0000000000000004_4572;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
  wire [31:0] _MUL826__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:972:131
  wire [31:0] _ADD825__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:971:130
  wire [31:0] _dup824__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:970:111
  wire [31:0] _dup824__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:970:111
  wire [31:0] _dup823__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:969:111
  wire [31:0] _dup823__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:969:111
  wire [31:0] _ADD822__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:968:130
  wire [31:0] _dup821_const_fix_32_0_1__0000000000002000_1950;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:967:473
  wire [31:0] _dup821_const_fix_32_0_1__0000000000002000_2314;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:967:473
  wire [31:0] _dup821_const_fix_32_0_1__0000000000002000_2678;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:967:473
  wire [31:0] _dup821_const_fix_32_0_1__0000000000002000_3042;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:967:473
  wire [31:0] _dup821_const_fix_32_0_1__0000000000002000_3406;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:967:473
  wire [31:0] _dup821_const_fix_32_0_1__0000000000002000_3770;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:967:473
  wire [31:0] _dup821_const_fix_32_0_1__0000000000002000_4134;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:967:473
  wire [31:0] _dup821_const_fix_32_0_1__0000000000002000_4498;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:967:473
  wire [31:0] _SHL8820__dfc_wire_1923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:966:89
  wire [31:0] _CAST819__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:965:84
  wire [31:0] _CAST818__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:964:84
  wire [31:0] _CAST817__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:963:84
  wire [31:0] _CAST816__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:962:84
  wire [31:0] _CAST815__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:961:84
  wire [31:0] _CAST814__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:960:84
  wire [31:0] _CAST813__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:959:84
  wire [31:0] _SHL8812__dfc_wire_1923;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:958:89
  wire [31:0] _CAST811__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:957:84
  wire [15:0] _CAST810__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:956:87
  wire [31:0] _SHR8809__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:955:87
  wire [31:0] _SUB808__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:954:109
  wire [15:0] _CAST807__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:953:87
  wire [31:0] _SHR8806__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:952:87
  wire [31:0] _SUB805__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:951:109
  wire [15:0] _CAST804__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:950:87
  wire [31:0] _SHR8803__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:949:87
  wire [31:0] _SUB802__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:948:109
  wire [15:0] _CAST801__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:947:87
  wire [31:0] _SHR8800__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:946:87
  wire [31:0] _SUB799__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:945:109
  wire [15:0] _CAST798__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:944:87
  wire [31:0] _SHR8797__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:943:87
  wire [31:0] _ADD796__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:942:130
  wire [31:0] _dup795__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:941:111
  wire [31:0] _dup795__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:941:111
  wire [31:0] _dup794__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:940:111
  wire [31:0] _dup794__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:940:111
  wire [15:0] _CAST793__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:939:87
  wire [31:0] _SHR8792__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:938:87
  wire [31:0] _ADD791__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:937:130
  wire [31:0] _dup790__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:936:111
  wire [31:0] _dup790__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:936:111
  wire [31:0] _dup789__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:935:111
  wire [31:0] _dup789__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:935:111
  wire [15:0] _CAST788__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:934:87
  wire [31:0] _SHR8787__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:933:87
  wire [31:0] _ADD786__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:932:130
  wire [31:0] _dup785__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:931:111
  wire [31:0] _dup785__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:931:111
  wire [31:0] _dup784__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:930:111
  wire [31:0] _dup784__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:930:111
  wire [15:0] _CAST783__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:929:87
  wire [31:0] _SHR8782__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:928:87
  wire [31:0] _ADD781__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:927:130
  wire [31:0] _dup780__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:926:111
  wire [31:0] _dup780__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:926:111
  wire [31:0] _dup779__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:925:111
  wire [31:0] _dup779__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:925:111
  wire [31:0] _SHR8778__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:924:87
  wire [31:0] _ADD777__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:923:130
  wire [31:0] _MUL776__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:922:131
  wire [31:0] _SUB775__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:921:109
  wire [31:0] _SHR8774__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:920:87
  wire [31:0] _ADD773__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:919:130
  wire [31:0] _MUL772__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:918:131
  wire [31:0] _ADD771__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:917:130
  wire [31:0] _dup770__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:916:111
  wire [31:0] _dup770__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:916:111
  wire [31:0] _dup769__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:915:111
  wire [31:0] _dup769__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:915:111
  wire [31:0] _SUB768__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:914:109
  wire [31:0] _ADD767__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:913:130
  wire [31:0] _dup766__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:912:111
  wire [31:0] _dup766__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:912:111
  wire [31:0] _dup765__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:911:111
  wire [31:0] _dup765__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:911:111
  wire [31:0] _SUB764__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:910:109
  wire [31:0] _ADD763__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:909:130
  wire [31:0] _dup762__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:908:111
  wire [31:0] _dup762__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:908:111
  wire [31:0] _dup761__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:907:111
  wire [31:0] _dup761__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:907:111
  wire [31:0] _SUB760__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:906:109
  wire [31:0] _ADD759__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:905:130
  wire [31:0] _dup758__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:904:111
  wire [31:0] _dup758__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:904:111
  wire [31:0] _dup757__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:903:111
  wire [31:0] _dup757__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:903:111
  wire [31:0] _SUB756__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:902:109
  wire [31:0] _ADD755__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:901:130
  wire [31:0] _dup754__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:900:111
  wire [31:0] _dup754__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:900:111
  wire [31:0] _dup753__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:899:111
  wire [31:0] _dup753__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:899:111
  wire [31:0] _ADD752__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:898:130
  wire [31:0] _MUL751__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:897:131
  wire [31:0] _SUB750__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:896:109
  wire [31:0] _dup749__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:895:111
  wire [31:0] _dup749__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:895:111
  wire [31:0] _MUL748__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:894:131
  wire [31:0] _MUL747__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:893:131
  wire [31:0] _ADD746__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:892:130
  wire [31:0] _dup745__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:891:111
  wire [31:0] _dup745__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:891:111
  wire [31:0] _dup744__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:890:111
  wire [31:0] _dup744__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:890:111
  wire [31:0] _SUB743__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:889:109
  wire [31:0] _ADD742__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:888:130
  wire [31:0] _dup741__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:887:111
  wire [31:0] _dup741__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:887:111
  wire [31:0] _dup740__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:886:111
  wire [31:0] _dup740__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:886:111
  wire [31:0] _SUB739__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:885:109
  wire [31:0] _MUL738__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:884:131
  wire [31:0] _SUB737__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:883:109
  wire [31:0] _dup736__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:882:111
  wire [31:0] _dup736__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:882:111
  wire [31:0] _MUL735__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:881:131
  wire [31:0] _MUL734__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:880:131
  wire [31:0] _ADD733__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:879:130
  wire [31:0] _dup732__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:878:111
  wire [31:0] _dup732__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:878:111
  wire [31:0] _dup731__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:877:111
  wire [31:0] _dup731__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:877:111
  wire [31:0] _SUB730__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:876:109
  wire [31:0] _MUL729__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:875:131
  wire [31:0] _ADD728__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:874:130
  wire [31:0] _dup727__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:873:111
  wire [31:0] _dup727__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:873:111
  wire [31:0] _MUL726__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:872:131
  wire [31:0] _MUL725__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:871:131
  wire [31:0] _ADD724__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:870:130
  wire [31:0] _dup723__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:869:111
  wire [31:0] _dup723__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:869:111
  wire [31:0] _dup722__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:868:111
  wire [31:0] _dup722__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:868:111
  wire [31:0] _ADD721__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:867:130
  wire [31:0] _SHL11720__dfc_wire_75;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:866:89
  wire [31:0] _CAST719__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:865:84
  wire [31:0] _CAST718__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:864:84
  wire [31:0] _CAST717__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:863:84
  wire [31:0] _CAST716__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:862:84
  wire [31:0] _CAST715__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:861:84
  wire [31:0] _CAST714__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:860:84
  wire [31:0] _CAST713__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:859:84
  wire [31:0] _SHL11712__dfc_wire_75;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:858:89
  wire [31:0] _CAST711__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:857:84
  wire [15:0] _CAST710__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:856:87
  wire [31:0] _SHR8709__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:855:87
  wire [31:0] _SUB708__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:854:109
  wire [15:0] _CAST707__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:853:87
  wire [31:0] _SHR8706__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:852:87
  wire [31:0] _SUB705__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:851:109
  wire [15:0] _CAST704__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:850:87
  wire [31:0] _SHR8703__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:849:87
  wire [31:0] _SUB702__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:848:109
  wire [15:0] _CAST701__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:847:87
  wire [31:0] _SHR8700__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:846:87
  wire [31:0] _SUB699__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:845:109
  wire [15:0] _CAST698__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:844:87
  wire [31:0] _SHR8697__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:843:87
  wire [31:0] _ADD696__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:842:130
  wire [31:0] _dup695__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:841:111
  wire [31:0] _dup695__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:841:111
  wire [31:0] _dup694__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:840:111
  wire [31:0] _dup694__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:840:111
  wire [15:0] _CAST693__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:839:87
  wire [31:0] _SHR8692__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:838:87
  wire [31:0] _ADD691__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:837:130
  wire [31:0] _dup690__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:836:111
  wire [31:0] _dup690__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:836:111
  wire [31:0] _dup689__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:835:111
  wire [31:0] _dup689__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:835:111
  wire [15:0] _CAST688__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:834:87
  wire [31:0] _SHR8687__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:833:87
  wire [31:0] _ADD686__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:832:130
  wire [31:0] _dup685__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:831:111
  wire [31:0] _dup685__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:831:111
  wire [31:0] _dup684__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:830:111
  wire [31:0] _dup684__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:830:111
  wire [15:0] _CAST683__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:829:87
  wire [31:0] _SHR8682__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:828:87
  wire [31:0] _ADD681__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:827:130
  wire [31:0] _dup680__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:826:111
  wire [31:0] _dup680__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:826:111
  wire [31:0] _dup679__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:825:111
  wire [31:0] _dup679__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:825:111
  wire [31:0] _SHR8678__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:824:87
  wire [31:0] _ADD677__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:823:130
  wire [31:0] _MUL676__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:822:131
  wire [31:0] _SUB675__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:821:109
  wire [31:0] _SHR8674__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:820:87
  wire [31:0] _ADD673__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:819:130
  wire [31:0] _MUL672__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:818:131
  wire [31:0] _ADD671__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:817:130
  wire [31:0] _dup670__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:816:111
  wire [31:0] _dup670__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:816:111
  wire [31:0] _dup669__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:815:111
  wire [31:0] _dup669__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:815:111
  wire [31:0] _SUB668__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:814:109
  wire [31:0] _ADD667__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:813:130
  wire [31:0] _dup666__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:812:111
  wire [31:0] _dup666__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:812:111
  wire [31:0] _dup665__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:811:111
  wire [31:0] _dup665__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:811:111
  wire [31:0] _SUB664__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:810:109
  wire [31:0] _ADD663__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:809:130
  wire [31:0] _dup662__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:808:111
  wire [31:0] _dup662__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:808:111
  wire [31:0] _dup661__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:807:111
  wire [31:0] _dup661__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:807:111
  wire [31:0] _SUB660__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:806:109
  wire [31:0] _ADD659__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:805:130
  wire [31:0] _dup658__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:804:111
  wire [31:0] _dup658__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:804:111
  wire [31:0] _dup657__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:803:111
  wire [31:0] _dup657__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:803:111
  wire [31:0] _SUB656__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:802:109
  wire [31:0] _ADD655__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:801:130
  wire [31:0] _dup654__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:800:111
  wire [31:0] _dup654__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:800:111
  wire [31:0] _dup653__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:799:111
  wire [31:0] _dup653__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:799:111
  wire [31:0] _ADD652__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:798:130
  wire [31:0] _MUL651__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:797:131
  wire [31:0] _SUB650__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:796:109
  wire [31:0] _dup649__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:795:111
  wire [31:0] _dup649__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:795:111
  wire [31:0] _MUL648__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:794:131
  wire [31:0] _MUL647__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:793:131
  wire [31:0] _ADD646__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:792:130
  wire [31:0] _dup645__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:791:111
  wire [31:0] _dup645__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:791:111
  wire [31:0] _dup644__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:790:111
  wire [31:0] _dup644__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:790:111
  wire [31:0] _SUB643__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:789:109
  wire [31:0] _ADD642__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:788:130
  wire [31:0] _dup641__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:787:111
  wire [31:0] _dup641__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:787:111
  wire [31:0] _dup640__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:786:111
  wire [31:0] _dup640__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:786:111
  wire [31:0] _SUB639__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:785:109
  wire [31:0] _MUL638__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:784:131
  wire [31:0] _SUB637__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:783:109
  wire [31:0] _dup636__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:782:111
  wire [31:0] _dup636__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:782:111
  wire [31:0] _MUL635__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:781:131
  wire [31:0] _MUL634__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:780:131
  wire [31:0] _ADD633__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:779:130
  wire [31:0] _dup632__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:778:111
  wire [31:0] _dup632__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:778:111
  wire [31:0] _dup631__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:777:111
  wire [31:0] _dup631__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:777:111
  wire [31:0] _SUB630__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:776:109
  wire [31:0] _MUL629__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:775:131
  wire [31:0] _ADD628__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:774:130
  wire [31:0] _dup627__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:773:111
  wire [31:0] _dup627__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:773:111
  wire [31:0] _MUL626__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:772:131
  wire [31:0] _MUL625__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:771:131
  wire [31:0] _ADD624__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:770:130
  wire [31:0] _dup623__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:769:111
  wire [31:0] _dup623__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:769:111
  wire [31:0] _dup622__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:768:111
  wire [31:0] _dup622__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:768:111
  wire [31:0] _ADD621__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:767:130
  wire [31:0] _SHL11620__dfc_wire_75;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:766:89
  wire [31:0] _CAST619__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:765:84
  wire [31:0] _CAST618__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:764:84
  wire [31:0] _CAST617__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:763:84
  wire [31:0] _CAST616__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:762:84
  wire [31:0] _CAST615__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:761:84
  wire [31:0] _CAST614__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:760:84
  wire [31:0] _CAST613__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:759:84
  wire [31:0] _SHL11612__dfc_wire_75;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:758:89
  wire [31:0] _CAST611__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:757:84
  wire [15:0] _CAST610__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:756:87
  wire [31:0] _SHR8609__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:755:87
  wire [31:0] _SUB608__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:754:109
  wire [15:0] _CAST607__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:753:87
  wire [31:0] _SHR8606__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:752:87
  wire [31:0] _SUB605__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:751:109
  wire [15:0] _CAST604__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:750:87
  wire [31:0] _SHR8603__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:749:87
  wire [31:0] _SUB602__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:748:109
  wire [15:0] _CAST601__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:747:87
  wire [31:0] _SHR8600__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:746:87
  wire [31:0] _SUB599__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:745:109
  wire [15:0] _CAST598__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:744:87
  wire [31:0] _SHR8597__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:743:87
  wire [31:0] _ADD596__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:742:130
  wire [31:0] _dup595__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:741:111
  wire [31:0] _dup595__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:741:111
  wire [31:0] _dup594__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:740:111
  wire [31:0] _dup594__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:740:111
  wire [15:0] _CAST593__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:739:87
  wire [31:0] _SHR8592__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:738:87
  wire [31:0] _ADD591__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:737:130
  wire [31:0] _dup590__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:736:111
  wire [31:0] _dup590__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:736:111
  wire [31:0] _dup589__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:735:111
  wire [31:0] _dup589__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:735:111
  wire [15:0] _CAST588__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:734:87
  wire [31:0] _SHR8587__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:733:87
  wire [31:0] _ADD586__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:732:130
  wire [31:0] _dup585__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:731:111
  wire [31:0] _dup585__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:731:111
  wire [31:0] _dup584__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:730:111
  wire [31:0] _dup584__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:730:111
  wire [15:0] _CAST583__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:729:87
  wire [31:0] _SHR8582__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:728:87
  wire [31:0] _ADD581__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:727:130
  wire [31:0] _dup580__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:726:111
  wire [31:0] _dup580__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:726:111
  wire [31:0] _dup579__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:725:111
  wire [31:0] _dup579__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:725:111
  wire [31:0] _SHR8578__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:724:87
  wire [31:0] _ADD577__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:723:130
  wire [31:0] _MUL576__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:722:131
  wire [31:0] _SUB575__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:721:109
  wire [31:0] _SHR8574__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:720:87
  wire [31:0] _ADD573__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:719:130
  wire [31:0] _MUL572__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:718:131
  wire [31:0] _ADD571__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:717:130
  wire [31:0] _dup570__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:716:111
  wire [31:0] _dup570__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:716:111
  wire [31:0] _dup569__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:715:111
  wire [31:0] _dup569__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:715:111
  wire [31:0] _SUB568__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:714:109
  wire [31:0] _ADD567__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:713:130
  wire [31:0] _dup566__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:712:111
  wire [31:0] _dup566__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:712:111
  wire [31:0] _dup565__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:711:111
  wire [31:0] _dup565__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:711:111
  wire [31:0] _SUB564__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:710:109
  wire [31:0] _ADD563__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:709:130
  wire [31:0] _dup562__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:708:111
  wire [31:0] _dup562__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:708:111
  wire [31:0] _dup561__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:707:111
  wire [31:0] _dup561__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:707:111
  wire [31:0] _SUB560__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:706:109
  wire [31:0] _ADD559__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:705:130
  wire [31:0] _dup558__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:704:111
  wire [31:0] _dup558__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:704:111
  wire [31:0] _dup557__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:703:111
  wire [31:0] _dup557__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:703:111
  wire [31:0] _SUB556__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:702:109
  wire [31:0] _ADD555__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:701:130
  wire [31:0] _dup554__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:700:111
  wire [31:0] _dup554__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:700:111
  wire [31:0] _dup553__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:699:111
  wire [31:0] _dup553__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:699:111
  wire [31:0] _ADD552__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:698:130
  wire [31:0] _MUL551__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:697:131
  wire [31:0] _SUB550__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:696:109
  wire [31:0] _dup549__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:695:111
  wire [31:0] _dup549__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:695:111
  wire [31:0] _MUL548__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:694:131
  wire [31:0] _MUL547__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:693:131
  wire [31:0] _ADD546__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:692:130
  wire [31:0] _dup545__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:691:111
  wire [31:0] _dup545__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:691:111
  wire [31:0] _dup544__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:690:111
  wire [31:0] _dup544__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:690:111
  wire [31:0] _SUB543__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:689:109
  wire [31:0] _ADD542__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:688:130
  wire [31:0] _dup541__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:687:111
  wire [31:0] _dup541__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:687:111
  wire [31:0] _dup540__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:686:111
  wire [31:0] _dup540__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:686:111
  wire [31:0] _SUB539__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:685:109
  wire [31:0] _MUL538__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:684:131
  wire [31:0] _SUB537__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:683:109
  wire [31:0] _dup536__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:682:111
  wire [31:0] _dup536__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:682:111
  wire [31:0] _MUL535__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:681:131
  wire [31:0] _MUL534__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:680:131
  wire [31:0] _ADD533__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:679:130
  wire [31:0] _dup532__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:678:111
  wire [31:0] _dup532__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:678:111
  wire [31:0] _dup531__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:677:111
  wire [31:0] _dup531__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:677:111
  wire [31:0] _SUB530__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:676:109
  wire [31:0] _MUL529__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:675:131
  wire [31:0] _ADD528__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:674:130
  wire [31:0] _dup527__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:673:111
  wire [31:0] _dup527__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:673:111
  wire [31:0] _MUL526__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:672:131
  wire [31:0] _MUL525__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:671:131
  wire [31:0] _ADD524__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:670:130
  wire [31:0] _dup523__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:669:111
  wire [31:0] _dup523__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:669:111
  wire [31:0] _dup522__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:668:111
  wire [31:0] _dup522__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:668:111
  wire [31:0] _ADD521__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:667:130
  wire [31:0] _SHL11520__dfc_wire_75;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:666:89
  wire [31:0] _CAST519__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:665:84
  wire [31:0] _CAST518__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:664:84
  wire [31:0] _CAST517__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:663:84
  wire [31:0] _CAST516__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:662:84
  wire [31:0] _CAST515__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:661:84
  wire [31:0] _CAST514__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:660:84
  wire [31:0] _CAST513__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:659:84
  wire [31:0] _SHL11512__dfc_wire_75;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:658:89
  wire [31:0] _CAST511__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:657:84
  wire [15:0] _CAST510__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:656:87
  wire [31:0] _SHR8509__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:655:87
  wire [31:0] _SUB508__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:654:109
  wire [15:0] _CAST507__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:653:87
  wire [31:0] _SHR8506__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:652:87
  wire [31:0] _SUB505__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:651:109
  wire [15:0] _CAST504__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:650:87
  wire [31:0] _SHR8503__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:649:87
  wire [31:0] _SUB502__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:648:109
  wire [15:0] _CAST501__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:647:87
  wire [31:0] _SHR8500__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:646:87
  wire [31:0] _SUB499__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:645:109
  wire [15:0] _CAST498__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:644:87
  wire [31:0] _SHR8497__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:643:87
  wire [31:0] _ADD496__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:642:130
  wire [31:0] _dup495__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:641:111
  wire [31:0] _dup495__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:641:111
  wire [31:0] _dup494__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:640:111
  wire [31:0] _dup494__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:640:111
  wire [15:0] _CAST493__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:639:87
  wire [31:0] _SHR8492__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:638:87
  wire [31:0] _ADD491__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:637:130
  wire [31:0] _dup490__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:636:111
  wire [31:0] _dup490__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:636:111
  wire [31:0] _dup489__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:635:111
  wire [31:0] _dup489__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:635:111
  wire [15:0] _CAST488__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:634:87
  wire [31:0] _SHR8487__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:633:87
  wire [31:0] _ADD486__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:632:130
  wire [31:0] _dup485__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:631:111
  wire [31:0] _dup485__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:631:111
  wire [31:0] _dup484__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:630:111
  wire [31:0] _dup484__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:630:111
  wire [15:0] _CAST483__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:629:87
  wire [31:0] _SHR8482__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:628:87
  wire [31:0] _ADD481__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:627:130
  wire [31:0] _dup480__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:626:111
  wire [31:0] _dup480__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:626:111
  wire [31:0] _dup479__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:625:111
  wire [31:0] _dup479__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:625:111
  wire [31:0] _SHR8478__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:624:87
  wire [31:0] _ADD477__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:623:130
  wire [31:0] _MUL476__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:622:131
  wire [31:0] _SUB475__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:621:109
  wire [31:0] _SHR8474__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:620:87
  wire [31:0] _ADD473__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:619:130
  wire [31:0] _MUL472__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:618:131
  wire [31:0] _ADD471__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:617:130
  wire [31:0] _dup470__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:616:111
  wire [31:0] _dup470__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:616:111
  wire [31:0] _dup469__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:615:111
  wire [31:0] _dup469__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:615:111
  wire [31:0] _SUB468__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:614:109
  wire [31:0] _ADD467__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:613:130
  wire [31:0] _dup466__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:612:111
  wire [31:0] _dup466__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:612:111
  wire [31:0] _dup465__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:611:111
  wire [31:0] _dup465__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:611:111
  wire [31:0] _SUB464__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:610:109
  wire [31:0] _ADD463__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:609:130
  wire [31:0] _dup462__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:608:111
  wire [31:0] _dup462__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:608:111
  wire [31:0] _dup461__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:607:111
  wire [31:0] _dup461__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:607:111
  wire [31:0] _SUB460__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:606:109
  wire [31:0] _ADD459__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:605:130
  wire [31:0] _dup458__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:604:111
  wire [31:0] _dup458__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:604:111
  wire [31:0] _dup457__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:603:111
  wire [31:0] _dup457__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:603:111
  wire [31:0] _SUB456__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:602:109
  wire [31:0] _ADD455__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:601:130
  wire [31:0] _dup454__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:600:111
  wire [31:0] _dup454__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:600:111
  wire [31:0] _dup453__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:599:111
  wire [31:0] _dup453__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:599:111
  wire [31:0] _ADD452__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:598:130
  wire [31:0] _MUL451__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:597:131
  wire [31:0] _SUB450__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:596:109
  wire [31:0] _dup449__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:595:111
  wire [31:0] _dup449__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:595:111
  wire [31:0] _MUL448__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:594:131
  wire [31:0] _MUL447__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:593:131
  wire [31:0] _ADD446__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:592:130
  wire [31:0] _dup445__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:591:111
  wire [31:0] _dup445__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:591:111
  wire [31:0] _dup444__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:590:111
  wire [31:0] _dup444__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:590:111
  wire [31:0] _SUB443__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:589:109
  wire [31:0] _ADD442__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:588:130
  wire [31:0] _dup441__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:587:111
  wire [31:0] _dup441__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:587:111
  wire [31:0] _dup440__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:586:111
  wire [31:0] _dup440__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:586:111
  wire [31:0] _SUB439__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:585:109
  wire [31:0] _MUL438__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:584:131
  wire [31:0] _SUB437__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:583:109
  wire [31:0] _dup436__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:582:111
  wire [31:0] _dup436__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:582:111
  wire [31:0] _MUL435__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:581:131
  wire [31:0] _MUL434__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:580:131
  wire [31:0] _ADD433__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:579:130
  wire [31:0] _dup432__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:578:111
  wire [31:0] _dup432__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:578:111
  wire [31:0] _dup431__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:577:111
  wire [31:0] _dup431__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:577:111
  wire [31:0] _SUB430__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:576:109
  wire [31:0] _MUL429__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:575:131
  wire [31:0] _ADD428__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:574:130
  wire [31:0] _dup427__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:573:111
  wire [31:0] _dup427__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:573:111
  wire [31:0] _MUL426__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:572:131
  wire [31:0] _MUL425__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:571:131
  wire [31:0] _ADD424__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:570:130
  wire [31:0] _dup423__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:569:111
  wire [31:0] _dup423__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:569:111
  wire [31:0] _dup422__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:568:111
  wire [31:0] _dup422__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:568:111
  wire [31:0] _ADD421__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:567:130
  wire [31:0] _SHL11420__dfc_wire_75;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:566:89
  wire [31:0] _CAST419__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:565:84
  wire [31:0] _CAST418__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:564:84
  wire [31:0] _CAST417__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:563:84
  wire [31:0] _CAST416__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:562:84
  wire [31:0] _CAST415__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:561:84
  wire [31:0] _CAST414__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:560:84
  wire [31:0] _CAST413__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:559:84
  wire [31:0] _SHL11412__dfc_wire_75;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:558:89
  wire [31:0] _CAST411__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:557:84
  wire [15:0] _CAST410__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:556:87
  wire [31:0] _SHR8409__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:555:87
  wire [31:0] _SUB408__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:554:109
  wire [15:0] _CAST407__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:553:87
  wire [31:0] _SHR8406__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:552:87
  wire [31:0] _SUB405__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:551:109
  wire [15:0] _CAST404__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:550:87
  wire [31:0] _SHR8403__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:549:87
  wire [31:0] _SUB402__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:548:109
  wire [15:0] _CAST401__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:547:87
  wire [31:0] _SHR8400__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:546:87
  wire [31:0] _SUB399__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:545:109
  wire [15:0] _CAST398__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:544:87
  wire [31:0] _SHR8397__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:543:87
  wire [31:0] _ADD396__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:542:130
  wire [31:0] _dup395__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:541:111
  wire [31:0] _dup395__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:541:111
  wire [31:0] _dup394__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:540:111
  wire [31:0] _dup394__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:540:111
  wire [15:0] _CAST393__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:539:87
  wire [31:0] _SHR8392__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:538:87
  wire [31:0] _ADD391__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:537:130
  wire [31:0] _dup390__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:536:111
  wire [31:0] _dup390__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:536:111
  wire [31:0] _dup389__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:535:111
  wire [31:0] _dup389__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:535:111
  wire [15:0] _CAST388__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:534:87
  wire [31:0] _SHR8387__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:533:87
  wire [31:0] _ADD386__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:532:130
  wire [31:0] _dup385__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:531:111
  wire [31:0] _dup385__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:531:111
  wire [31:0] _dup384__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:530:111
  wire [31:0] _dup384__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:530:111
  wire [15:0] _CAST383__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:529:87
  wire [31:0] _SHR8382__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:528:87
  wire [31:0] _ADD381__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:527:130
  wire [31:0] _dup380__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:526:111
  wire [31:0] _dup380__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:526:111
  wire [31:0] _dup379__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:525:111
  wire [31:0] _dup379__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:525:111
  wire [31:0] _SHR8378__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:524:87
  wire [31:0] _ADD377__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:523:130
  wire [31:0] _MUL376__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:522:131
  wire [31:0] _SUB375__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:521:109
  wire [31:0] _SHR8374__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:520:87
  wire [31:0] _ADD373__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:519:130
  wire [31:0] _MUL372__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:518:131
  wire [31:0] _ADD371__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:517:130
  wire [31:0] _dup370__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:516:111
  wire [31:0] _dup370__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:516:111
  wire [31:0] _dup369__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:515:111
  wire [31:0] _dup369__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:515:111
  wire [31:0] _SUB368__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:514:109
  wire [31:0] _ADD367__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:513:130
  wire [31:0] _dup366__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:512:111
  wire [31:0] _dup366__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:512:111
  wire [31:0] _dup365__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:511:111
  wire [31:0] _dup365__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:511:111
  wire [31:0] _SUB364__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:510:109
  wire [31:0] _ADD363__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:509:130
  wire [31:0] _dup362__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:508:111
  wire [31:0] _dup362__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:508:111
  wire [31:0] _dup361__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:507:111
  wire [31:0] _dup361__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:507:111
  wire [31:0] _SUB360__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:506:109
  wire [31:0] _ADD359__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:505:130
  wire [31:0] _dup358__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:504:111
  wire [31:0] _dup358__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:504:111
  wire [31:0] _dup357__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:503:111
  wire [31:0] _dup357__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:503:111
  wire [31:0] _SUB356__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:502:109
  wire [31:0] _ADD355__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:501:130
  wire [31:0] _dup354__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:500:111
  wire [31:0] _dup354__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:500:111
  wire [31:0] _dup353__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:499:111
  wire [31:0] _dup353__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:499:111
  wire [31:0] _ADD352__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:498:130
  wire [31:0] _MUL351__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:497:131
  wire [31:0] _SUB350__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:496:109
  wire [31:0] _dup349__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:495:111
  wire [31:0] _dup349__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:495:111
  wire [31:0] _MUL348__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:494:131
  wire [31:0] _MUL347__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:493:131
  wire [31:0] _ADD346__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:492:130
  wire [31:0] _dup345__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:491:111
  wire [31:0] _dup345__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:491:111
  wire [31:0] _dup344__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:490:111
  wire [31:0] _dup344__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:490:111
  wire [31:0] _SUB343__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:489:109
  wire [31:0] _ADD342__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:488:130
  wire [31:0] _dup341__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:487:111
  wire [31:0] _dup341__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:487:111
  wire [31:0] _dup340__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:486:111
  wire [31:0] _dup340__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:486:111
  wire [31:0] _SUB339__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:485:109
  wire [31:0] _MUL338__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:484:131
  wire [31:0] _SUB337__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:483:109
  wire [31:0] _dup336__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:482:111
  wire [31:0] _dup336__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:482:111
  wire [31:0] _MUL335__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:481:131
  wire [31:0] _MUL334__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:480:131
  wire [31:0] _ADD333__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:479:130
  wire [31:0] _dup332__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:478:111
  wire [31:0] _dup332__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:478:111
  wire [31:0] _dup331__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:477:111
  wire [31:0] _dup331__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:477:111
  wire [31:0] _SUB330__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:476:109
  wire [31:0] _MUL329__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:475:131
  wire [31:0] _ADD328__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:474:130
  wire [31:0] _dup327__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:473:111
  wire [31:0] _dup327__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:473:111
  wire [31:0] _MUL326__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:472:131
  wire [31:0] _MUL325__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:471:131
  wire [31:0] _ADD324__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:470:130
  wire [31:0] _dup323__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:469:111
  wire [31:0] _dup323__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:469:111
  wire [31:0] _dup322__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:468:111
  wire [31:0] _dup322__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:468:111
  wire [31:0] _ADD321__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:467:130
  wire [31:0] _SHL11320__dfc_wire_75;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:466:89
  wire [31:0] _CAST319__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:465:84
  wire [31:0] _CAST318__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:464:84
  wire [31:0] _CAST317__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:463:84
  wire [31:0] _CAST316__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:462:84
  wire [31:0] _CAST315__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:461:84
  wire [31:0] _CAST314__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:460:84
  wire [31:0] _CAST313__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:459:84
  wire [31:0] _SHL11312__dfc_wire_75;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:458:89
  wire [31:0] _CAST311__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:457:84
  wire [15:0] _CAST310__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:456:87
  wire [31:0] _SHR8309__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:455:87
  wire [31:0] _SUB308__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:454:109
  wire [15:0] _CAST307__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:453:87
  wire [31:0] _SHR8306__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:452:87
  wire [31:0] _SUB305__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:451:109
  wire [15:0] _CAST304__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:450:87
  wire [31:0] _SHR8303__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:449:87
  wire [31:0] _SUB302__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:448:109
  wire [15:0] _CAST301__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:447:87
  wire [31:0] _SHR8300__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:446:87
  wire [31:0] _SUB299__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:445:109
  wire [15:0] _CAST298__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:444:87
  wire [31:0] _SHR8297__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:443:87
  wire [31:0] _ADD296__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:442:130
  wire [31:0] _dup295__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:441:111
  wire [31:0] _dup295__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:441:111
  wire [31:0] _dup294__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:440:111
  wire [31:0] _dup294__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:440:111
  wire [15:0] _CAST293__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:439:87
  wire [31:0] _SHR8292__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:438:87
  wire [31:0] _ADD291__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:437:130
  wire [31:0] _dup290__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:436:111
  wire [31:0] _dup290__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:436:111
  wire [31:0] _dup289__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:435:111
  wire [31:0] _dup289__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:435:111
  wire [15:0] _CAST288__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:434:87
  wire [31:0] _SHR8287__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:433:87
  wire [31:0] _ADD286__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:432:130
  wire [31:0] _dup285__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:431:111
  wire [31:0] _dup285__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:431:111
  wire [31:0] _dup284__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:430:111
  wire [31:0] _dup284__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:430:111
  wire [15:0] _CAST283__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:429:87
  wire [31:0] _SHR8282__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:428:87
  wire [31:0] _ADD281__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:427:130
  wire [31:0] _dup280__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:426:111
  wire [31:0] _dup280__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:426:111
  wire [31:0] _dup279__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:425:111
  wire [31:0] _dup279__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:425:111
  wire [31:0] _SHR8278__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:424:87
  wire [31:0] _ADD277__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:423:130
  wire [31:0] _MUL276__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:422:131
  wire [31:0] _SUB275__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:421:109
  wire [31:0] _SHR8274__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:420:87
  wire [31:0] _ADD273__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:419:130
  wire [31:0] _MUL272__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:418:131
  wire [31:0] _ADD271__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:417:130
  wire [31:0] _dup270__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:416:111
  wire [31:0] _dup270__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:416:111
  wire [31:0] _dup269__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:415:111
  wire [31:0] _dup269__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:415:111
  wire [31:0] _SUB268__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:414:109
  wire [31:0] _ADD267__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:413:130
  wire [31:0] _dup266__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:412:111
  wire [31:0] _dup266__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:412:111
  wire [31:0] _dup265__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:411:111
  wire [31:0] _dup265__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:411:111
  wire [31:0] _SUB264__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:410:109
  wire [31:0] _ADD263__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:409:130
  wire [31:0] _dup262__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:408:111
  wire [31:0] _dup262__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:408:111
  wire [31:0] _dup261__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:407:111
  wire [31:0] _dup261__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:407:111
  wire [31:0] _SUB260__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:406:109
  wire [31:0] _ADD259__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:405:130
  wire [31:0] _dup258__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:404:111
  wire [31:0] _dup258__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:404:111
  wire [31:0] _dup257__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:403:111
  wire [31:0] _dup257__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:403:111
  wire [31:0] _SUB256__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:402:109
  wire [31:0] _ADD255__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:401:130
  wire [31:0] _dup254__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:400:111
  wire [31:0] _dup254__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:400:111
  wire [31:0] _dup253__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:399:111
  wire [31:0] _dup253__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:399:111
  wire [31:0] _ADD252__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:398:130
  wire [31:0] _MUL251__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:397:131
  wire [31:0] _SUB250__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:396:109
  wire [31:0] _dup249__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:395:111
  wire [31:0] _dup249__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:395:111
  wire [31:0] _MUL248__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:394:131
  wire [31:0] _MUL247__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:393:131
  wire [31:0] _ADD246__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:392:130
  wire [31:0] _dup245__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:391:111
  wire [31:0] _dup245__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:391:111
  wire [31:0] _dup244__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:390:111
  wire [31:0] _dup244__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:390:111
  wire [31:0] _SUB243__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:389:109
  wire [31:0] _ADD242__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:388:130
  wire [31:0] _dup241__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:387:111
  wire [31:0] _dup241__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:387:111
  wire [31:0] _dup240__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:386:111
  wire [31:0] _dup240__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:386:111
  wire [31:0] _SUB239__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:385:109
  wire [31:0] _MUL238__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:384:131
  wire [31:0] _SUB237__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:383:109
  wire [31:0] _dup236__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:382:111
  wire [31:0] _dup236__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:382:111
  wire [31:0] _MUL235__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:381:131
  wire [31:0] _MUL234__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:380:131
  wire [31:0] _ADD233__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:379:130
  wire [31:0] _dup232__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:378:111
  wire [31:0] _dup232__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:378:111
  wire [31:0] _dup231__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:377:111
  wire [31:0] _dup231__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:377:111
  wire [31:0] _SUB230__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:376:109
  wire [31:0] _MUL229__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:375:131
  wire [31:0] _ADD228__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:374:130
  wire [31:0] _dup227__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:373:111
  wire [31:0] _dup227__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:373:111
  wire [31:0] _MUL226__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:372:131
  wire [31:0] _MUL225__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:371:131
  wire [31:0] _ADD224__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:370:130
  wire [31:0] _dup223__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:369:111
  wire [31:0] _dup223__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:369:111
  wire [31:0] _dup222__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:368:111
  wire [31:0] _dup222__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:368:111
  wire [31:0] _ADD221__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:367:130
  wire [31:0] _SHL11220__dfc_wire_75;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:366:89
  wire [31:0] _CAST219__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:365:84
  wire [31:0] _CAST218__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:364:84
  wire [31:0] _CAST217__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:363:84
  wire [31:0] _CAST216__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:362:84
  wire [31:0] _CAST215__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:361:84
  wire [31:0] _CAST214__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:360:84
  wire [31:0] _CAST213__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:359:84
  wire [31:0] _SHL11212__dfc_wire_75;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:358:89
  wire [31:0] _CAST211__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:357:84
  wire [15:0] _CAST210__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:356:87
  wire [31:0] _SHR8209__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:355:87
  wire [31:0] _SUB208__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:354:109
  wire [15:0] _CAST207__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:353:87
  wire [31:0] _SHR8206__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:352:87
  wire [31:0] _SUB205__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:351:109
  wire [15:0] _CAST204__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:350:87
  wire [31:0] _SHR8203__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:349:87
  wire [31:0] _SUB202__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:348:109
  wire [15:0] _CAST201__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:347:87
  wire [31:0] _SHR8200__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:346:87
  wire [31:0] _SUB199__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:345:109
  wire [15:0] _CAST198__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:344:87
  wire [31:0] _SHR8197__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:343:87
  wire [31:0] _ADD196__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:342:130
  wire [31:0] _dup195__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:341:111
  wire [31:0] _dup195__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:341:111
  wire [31:0] _dup194__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:340:111
  wire [31:0] _dup194__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:340:111
  wire [15:0] _CAST193__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:339:87
  wire [31:0] _SHR8192__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:338:87
  wire [31:0] _ADD191__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:337:130
  wire [31:0] _dup190__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:336:111
  wire [31:0] _dup190__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:336:111
  wire [31:0] _dup189__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:335:111
  wire [31:0] _dup189__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:335:111
  wire [15:0] _CAST188__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:334:87
  wire [31:0] _SHR8187__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:333:87
  wire [31:0] _ADD186__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:332:130
  wire [31:0] _dup185__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:331:111
  wire [31:0] _dup185__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:331:111
  wire [31:0] _dup184__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:330:111
  wire [31:0] _dup184__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:330:111
  wire [15:0] _CAST183__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:329:87
  wire [31:0] _SHR8182__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:328:87
  wire [31:0] _ADD181__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:327:130
  wire [31:0] _dup180__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:326:111
  wire [31:0] _dup180__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:326:111
  wire [31:0] _dup179__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:325:111
  wire [31:0] _dup179__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:325:111
  wire [31:0] _SHR8178__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:324:87
  wire [31:0] _ADD177__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:323:130
  wire [31:0] _MUL176__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:322:131
  wire [31:0] _SUB175__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:321:109
  wire [31:0] _SHR8174__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:320:87
  wire [31:0] _ADD173__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:319:130
  wire [31:0] _MUL172__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:318:131
  wire [31:0] _ADD171__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:317:130
  wire [31:0] _dup170__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:316:111
  wire [31:0] _dup170__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:316:111
  wire [31:0] _dup169__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:315:111
  wire [31:0] _dup169__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:315:111
  wire [31:0] _SUB168__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:314:109
  wire [31:0] _ADD167__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:313:130
  wire [31:0] _dup166__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:312:111
  wire [31:0] _dup166__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:312:111
  wire [31:0] _dup165__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:311:111
  wire [31:0] _dup165__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:311:111
  wire [31:0] _SUB164__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:310:109
  wire [31:0] _ADD163__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:309:130
  wire [31:0] _dup162__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:308:111
  wire [31:0] _dup162__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:308:111
  wire [31:0] _dup161__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:307:111
  wire [31:0] _dup161__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:307:111
  wire [31:0] _SUB160__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:306:109
  wire [31:0] _ADD159__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:305:130
  wire [31:0] _dup158__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:304:111
  wire [31:0] _dup158__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:304:111
  wire [31:0] _dup157__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:303:111
  wire [31:0] _dup157__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:303:111
  wire [31:0] _SUB156__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:302:109
  wire [31:0] _ADD155__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:301:130
  wire [31:0] _dup154__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:300:111
  wire [31:0] _dup154__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:300:111
  wire [31:0] _dup153__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:299:111
  wire [31:0] _dup153__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:299:111
  wire [31:0] _ADD152__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:298:130
  wire [31:0] _MUL151__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:297:131
  wire [31:0] _SUB150__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:296:109
  wire [31:0] _dup149__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:295:111
  wire [31:0] _dup149__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:295:111
  wire [31:0] _MUL148__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:294:131
  wire [31:0] _MUL147__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:293:131
  wire [31:0] _ADD146__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:292:130
  wire [31:0] _dup145__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:291:111
  wire [31:0] _dup145__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:291:111
  wire [31:0] _dup144__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:290:111
  wire [31:0] _dup144__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:290:111
  wire [31:0] _SUB143__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:289:109
  wire [31:0] _ADD142__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:288:130
  wire [31:0] _dup141__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:287:111
  wire [31:0] _dup141__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:287:111
  wire [31:0] _dup140__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:286:111
  wire [31:0] _dup140__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:286:111
  wire [31:0] _SUB139__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:285:109
  wire [31:0] _MUL138__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:284:131
  wire [31:0] _SUB137__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:283:109
  wire [31:0] _dup136__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:282:111
  wire [31:0] _dup136__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:282:111
  wire [31:0] _MUL135__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:281:131
  wire [31:0] _MUL134__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:280:131
  wire [31:0] _ADD133__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:279:130
  wire [31:0] _dup132__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:278:111
  wire [31:0] _dup132__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:278:111
  wire [31:0] _dup131__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:277:111
  wire [31:0] _dup131__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:277:111
  wire [31:0] _SUB130__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:276:109
  wire [31:0] _MUL129__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:275:131
  wire [31:0] _ADD128__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:274:130
  wire [31:0] _dup127__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:273:111
  wire [31:0] _dup127__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:273:111
  wire [31:0] _MUL126__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:272:131
  wire [31:0] _MUL125__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:271:131
  wire [31:0] _ADD124__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:270:130
  wire [31:0] _dup123__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:269:111
  wire [31:0] _dup123__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:269:111
  wire [31:0] _dup122__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:268:111
  wire [31:0] _dup122__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:268:111
  wire [31:0] _ADD121__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:267:130
  wire [31:0] _SHL11120__dfc_wire_75;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:266:89
  wire [31:0] _CAST119__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:265:84
  wire [31:0] _CAST118__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:264:84
  wire [31:0] _CAST117__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:263:84
  wire [31:0] _CAST116__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:262:84
  wire [31:0] _CAST115__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:261:84
  wire [31:0] _CAST114__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:260:84
  wire [31:0] _CAST113__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:259:84
  wire [31:0] _SHL11112__dfc_wire_75;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:258:89
  wire [31:0] _CAST111__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:257:84
  wire [15:0] _CAST110__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:256:87
  wire [31:0] _SHR8109__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:255:87
  wire [31:0] _SUB108__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:254:109
  wire [15:0] _CAST107__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:253:87
  wire [31:0] _SHR8106__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:252:87
  wire [31:0] _SUB105__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:251:109
  wire [15:0] _CAST104__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:250:87
  wire [31:0] _SHR8103__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:249:87
  wire [31:0] _SUB102__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:248:109
  wire [15:0] _CAST101__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:247:87
  wire [31:0] _SHR8100__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:246:87
  wire [31:0] _SUB99__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:245:104
  wire [15:0] _CAST98__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:244:83
  wire [31:0] _SHR897__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:243:83
  wire [31:0] _ADD96__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:242:125
  wire [31:0] _dup95__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:241:106
  wire [31:0] _dup95__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:241:106
  wire [31:0] _dup94__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:240:106
  wire [31:0] _dup94__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:240:106
  wire [15:0] _CAST93__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:239:83
  wire [31:0] _SHR892__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:238:83
  wire [31:0] _ADD91__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:237:125
  wire [31:0] _dup90__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:236:106
  wire [31:0] _dup90__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:236:106
  wire [31:0] _dup89__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:235:106
  wire [31:0] _dup89__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:235:106
  wire [15:0] _CAST88__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:234:83
  wire [31:0] _SHR887__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:233:83
  wire [31:0] _ADD86__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:232:125
  wire [31:0] _dup85__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:231:106
  wire [31:0] _dup85__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:231:106
  wire [31:0] _dup84__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:230:106
  wire [31:0] _dup84__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:230:106
  wire [15:0] _CAST83__dfc_wire_236;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:229:83
  wire [31:0] _SHR882__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:228:83
  wire [31:0] _ADD81__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:227:125
  wire [31:0] _dup80__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:226:106
  wire [31:0] _dup80__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:226:106
  wire [31:0] _dup79__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:225:106
  wire [31:0] _dup79__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:225:106
  wire [31:0] _SHR878__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:224:83
  wire [31:0] _ADD77__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:223:125
  wire [31:0] _MUL76__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:222:126
  wire [31:0] _SUB75__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:221:104
  wire [31:0] _SHR874__dfc_wire_216;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:220:83
  wire [31:0] _ADD73__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:219:125
  wire [31:0] _MUL72__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:218:126
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_211;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_223;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_442;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_454;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_673;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_685;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_904;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_916;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_1135;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_1147;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_1366;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_1378;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_1597;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_1609;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_1828;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_1840;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_2080;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_2092;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_2444;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_2456;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_2808;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_2820;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_3172;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_3184;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_3536;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_3548;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_3900;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_3912;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_4264;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_4276;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_4628;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _dup71_const_fix_32_0_1__00000000000000b5_4640;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
  wire [31:0] _ADD70__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:216:125
  wire [31:0] _dup69__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:215:106
  wire [31:0] _dup69__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:215:106
  wire [31:0] _dup68__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:214:106
  wire [31:0] _dup68__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:214:106
  wire [31:0] _SUB67__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:213:104
  wire [31:0] _ADD66__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:212:125
  wire [31:0] _dup65__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:211:106
  wire [31:0] _dup65__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:211:106
  wire [31:0] _dup64__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:210:106
  wire [31:0] _dup64__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:210:106
  wire [31:0] _SUB63__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:209:104
  wire [31:0] _ADD62__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:208:125
  wire [31:0] _dup61__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:207:106
  wire [31:0] _dup61__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:207:106
  wire [31:0] _dup60__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:206:106
  wire [31:0] _dup60__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:206:106
  wire [31:0] _SUB59__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:205:104
  wire [31:0] _ADD58__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:204:125
  wire [31:0] _dup57__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:203:106
  wire [31:0] _dup57__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:203:106
  wire [31:0] _dup56__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:202:106
  wire [31:0] _dup56__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:202:106
  wire [31:0] _SUB55__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:201:104
  wire [31:0] _ADD54__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:200:125
  wire [31:0] _dup53__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:199:106
  wire [31:0] _dup53__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:199:106
  wire [31:0] _dup52__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:198:106
  wire [31:0] _dup52__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:198:106
  wire [31:0] _ADD51__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:197:125
  wire [31:0] _MUL50__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:196:126
  wire [31:0] _dup49_const_fix_32_0_1__0000000000000235_108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
  wire [31:0] _dup49_const_fix_32_0_1__0000000000000235_339;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
  wire [31:0] _dup49_const_fix_32_0_1__0000000000000235_570;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
  wire [31:0] _dup49_const_fix_32_0_1__0000000000000235_801;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
  wire [31:0] _dup49_const_fix_32_0_1__0000000000000235_1032;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
  wire [31:0] _dup49_const_fix_32_0_1__0000000000000235_1263;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
  wire [31:0] _dup49_const_fix_32_0_1__0000000000000235_1494;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
  wire [31:0] _dup49_const_fix_32_0_1__0000000000000235_1725;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
  wire [31:0] _dup49_const_fix_32_0_1__0000000000000235_1956;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
  wire [31:0] _dup49_const_fix_32_0_1__0000000000000235_2320;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
  wire [31:0] _dup49_const_fix_32_0_1__0000000000000235_2684;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
  wire [31:0] _dup49_const_fix_32_0_1__0000000000000235_3048;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
  wire [31:0] _dup49_const_fix_32_0_1__0000000000000235_3412;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
  wire [31:0] _dup49_const_fix_32_0_1__0000000000000235_3776;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
  wire [31:0] _dup49_const_fix_32_0_1__0000000000000235_4140;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
  wire [31:0] _dup49_const_fix_32_0_1__0000000000000235_4504;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
  wire [31:0] _SUB48__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:194:104
  wire [31:0] _dup47__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:193:106
  wire [31:0] _dup47__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:193:106
  wire [31:0] _MUL46__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:192:126
  wire [31:0] _dup45_const_fix_32_0_1__0000000000000235_108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
  wire [31:0] _dup45_const_fix_32_0_1__0000000000000235_339;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
  wire [31:0] _dup45_const_fix_32_0_1__0000000000000235_570;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
  wire [31:0] _dup45_const_fix_32_0_1__0000000000000235_801;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
  wire [31:0] _dup45_const_fix_32_0_1__0000000000000235_1032;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
  wire [31:0] _dup45_const_fix_32_0_1__0000000000000235_1263;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
  wire [31:0] _dup45_const_fix_32_0_1__0000000000000235_1494;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
  wire [31:0] _dup45_const_fix_32_0_1__0000000000000235_1725;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
  wire [31:0] _dup45_const_fix_32_0_1__0000000000000235_1956;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
  wire [31:0] _dup45_const_fix_32_0_1__0000000000000235_2320;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
  wire [31:0] _dup45_const_fix_32_0_1__0000000000000235_2684;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
  wire [31:0] _dup45_const_fix_32_0_1__0000000000000235_3048;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
  wire [31:0] _dup45_const_fix_32_0_1__0000000000000235_3412;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
  wire [31:0] _dup45_const_fix_32_0_1__0000000000000235_3776;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
  wire [31:0] _dup45_const_fix_32_0_1__0000000000000235_4140;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
  wire [31:0] _dup45_const_fix_32_0_1__0000000000000235_4504;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
  wire [31:0] _MUL44__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:190:126
  wire [31:0] _dup43_const_fix_32_0_1__0000000000000235_108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
  wire [31:0] _dup43_const_fix_32_0_1__0000000000000235_339;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
  wire [31:0] _dup43_const_fix_32_0_1__0000000000000235_570;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
  wire [31:0] _dup43_const_fix_32_0_1__0000000000000235_801;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
  wire [31:0] _dup43_const_fix_32_0_1__0000000000000235_1032;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
  wire [31:0] _dup43_const_fix_32_0_1__0000000000000235_1263;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
  wire [31:0] _dup43_const_fix_32_0_1__0000000000000235_1494;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
  wire [31:0] _dup43_const_fix_32_0_1__0000000000000235_1725;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
  wire [31:0] _dup43_const_fix_32_0_1__0000000000000235_1956;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
  wire [31:0] _dup43_const_fix_32_0_1__0000000000000235_2320;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
  wire [31:0] _dup43_const_fix_32_0_1__0000000000000235_2684;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
  wire [31:0] _dup43_const_fix_32_0_1__0000000000000235_3048;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
  wire [31:0] _dup43_const_fix_32_0_1__0000000000000235_3412;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
  wire [31:0] _dup43_const_fix_32_0_1__0000000000000235_3776;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
  wire [31:0] _dup43_const_fix_32_0_1__0000000000000235_4140;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
  wire [31:0] _dup43_const_fix_32_0_1__0000000000000235_4504;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
  wire [31:0] _ADD42__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:188:125
  wire [31:0] _dup41__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:187:106
  wire [31:0] _dup41__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:187:106
  wire [31:0] _dup40__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:186:106
  wire [31:0] _dup40__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:186:106
  wire [31:0] _SUB39__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:185:104
  wire [31:0] _ADD38__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:184:125
  wire [31:0] _dup37__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:183:106
  wire [31:0] _dup37__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:183:106
  wire [31:0] _dup36__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:182:106
  wire [31:0] _dup36__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:182:106
  wire [31:0] _SUB35__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:181:104
  wire [31:0] _MUL34__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:180:126
  wire [31:0] _dup33_const_fix_32_0_1__0000000000000235_108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
  wire [31:0] _dup33_const_fix_32_0_1__0000000000000235_339;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
  wire [31:0] _dup33_const_fix_32_0_1__0000000000000235_570;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
  wire [31:0] _dup33_const_fix_32_0_1__0000000000000235_801;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
  wire [31:0] _dup33_const_fix_32_0_1__0000000000000235_1032;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
  wire [31:0] _dup33_const_fix_32_0_1__0000000000000235_1263;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
  wire [31:0] _dup33_const_fix_32_0_1__0000000000000235_1494;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
  wire [31:0] _dup33_const_fix_32_0_1__0000000000000235_1725;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
  wire [31:0] _dup33_const_fix_32_0_1__0000000000000235_1956;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
  wire [31:0] _dup33_const_fix_32_0_1__0000000000000235_2320;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
  wire [31:0] _dup33_const_fix_32_0_1__0000000000000235_2684;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
  wire [31:0] _dup33_const_fix_32_0_1__0000000000000235_3048;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
  wire [31:0] _dup33_const_fix_32_0_1__0000000000000235_3412;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
  wire [31:0] _dup33_const_fix_32_0_1__0000000000000235_3776;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
  wire [31:0] _dup33_const_fix_32_0_1__0000000000000235_4140;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
  wire [31:0] _dup33_const_fix_32_0_1__0000000000000235_4504;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
  wire [31:0] _SUB32__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:178:104
  wire [31:0] _dup31__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:177:106
  wire [31:0] _dup31__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:177:106
  wire [31:0] _MUL30__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:176:126
  wire [31:0] _dup29_const_fix_32_0_1__0000000000000235_108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
  wire [31:0] _dup29_const_fix_32_0_1__0000000000000235_339;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
  wire [31:0] _dup29_const_fix_32_0_1__0000000000000235_570;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
  wire [31:0] _dup29_const_fix_32_0_1__0000000000000235_801;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
  wire [31:0] _dup29_const_fix_32_0_1__0000000000000235_1032;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
  wire [31:0] _dup29_const_fix_32_0_1__0000000000000235_1263;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
  wire [31:0] _dup29_const_fix_32_0_1__0000000000000235_1494;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
  wire [31:0] _dup29_const_fix_32_0_1__0000000000000235_1725;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
  wire [31:0] _dup29_const_fix_32_0_1__0000000000000235_1956;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
  wire [31:0] _dup29_const_fix_32_0_1__0000000000000235_2320;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
  wire [31:0] _dup29_const_fix_32_0_1__0000000000000235_2684;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
  wire [31:0] _dup29_const_fix_32_0_1__0000000000000235_3048;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
  wire [31:0] _dup29_const_fix_32_0_1__0000000000000235_3412;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
  wire [31:0] _dup29_const_fix_32_0_1__0000000000000235_3776;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
  wire [31:0] _dup29_const_fix_32_0_1__0000000000000235_4140;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
  wire [31:0] _dup29_const_fix_32_0_1__0000000000000235_4504;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
  wire [31:0] _MUL28__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:174:126
  wire [31:0] _dup27_const_fix_32_0_1__0000000000000235_108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
  wire [31:0] _dup27_const_fix_32_0_1__0000000000000235_339;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
  wire [31:0] _dup27_const_fix_32_0_1__0000000000000235_570;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
  wire [31:0] _dup27_const_fix_32_0_1__0000000000000235_801;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
  wire [31:0] _dup27_const_fix_32_0_1__0000000000000235_1032;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
  wire [31:0] _dup27_const_fix_32_0_1__0000000000000235_1263;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
  wire [31:0] _dup27_const_fix_32_0_1__0000000000000235_1494;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
  wire [31:0] _dup27_const_fix_32_0_1__0000000000000235_1725;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
  wire [31:0] _dup27_const_fix_32_0_1__0000000000000235_1956;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
  wire [31:0] _dup27_const_fix_32_0_1__0000000000000235_2320;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
  wire [31:0] _dup27_const_fix_32_0_1__0000000000000235_2684;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
  wire [31:0] _dup27_const_fix_32_0_1__0000000000000235_3048;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
  wire [31:0] _dup27_const_fix_32_0_1__0000000000000235_3412;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
  wire [31:0] _dup27_const_fix_32_0_1__0000000000000235_3776;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
  wire [31:0] _dup27_const_fix_32_0_1__0000000000000235_4140;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
  wire [31:0] _dup27_const_fix_32_0_1__0000000000000235_4504;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
  wire [31:0] _ADD26__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:172:125
  wire [31:0] _dup25__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:171:106
  wire [31:0] _dup25__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:171:106
  wire [31:0] _dup24__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:170:106
  wire [31:0] _dup24__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:170:106
  wire [31:0] _SUB23__dfc_wire_121;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:169:104
  wire [31:0] _MUL22__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:168:126
  wire [31:0] _dup21_const_fix_32_0_1__0000000000000235_108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
  wire [31:0] _dup21_const_fix_32_0_1__0000000000000235_339;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
  wire [31:0] _dup21_const_fix_32_0_1__0000000000000235_570;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
  wire [31:0] _dup21_const_fix_32_0_1__0000000000000235_801;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
  wire [31:0] _dup21_const_fix_32_0_1__0000000000000235_1032;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
  wire [31:0] _dup21_const_fix_32_0_1__0000000000000235_1263;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
  wire [31:0] _dup21_const_fix_32_0_1__0000000000000235_1494;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
  wire [31:0] _dup21_const_fix_32_0_1__0000000000000235_1725;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
  wire [31:0] _dup21_const_fix_32_0_1__0000000000000235_1956;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
  wire [31:0] _dup21_const_fix_32_0_1__0000000000000235_2320;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
  wire [31:0] _dup21_const_fix_32_0_1__0000000000000235_2684;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
  wire [31:0] _dup21_const_fix_32_0_1__0000000000000235_3048;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
  wire [31:0] _dup21_const_fix_32_0_1__0000000000000235_3412;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
  wire [31:0] _dup21_const_fix_32_0_1__0000000000000235_3776;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
  wire [31:0] _dup21_const_fix_32_0_1__0000000000000235_4140;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
  wire [31:0] _dup21_const_fix_32_0_1__0000000000000235_4504;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
  wire [31:0] _ADD20__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:166:125
  wire [31:0] _dup19__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:165:106
  wire [31:0] _dup19__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:165:106
  wire [31:0] _MUL18__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:164:126
  wire [31:0] _dup17_const_fix_32_0_1__0000000000000235_108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
  wire [31:0] _dup17_const_fix_32_0_1__0000000000000235_339;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
  wire [31:0] _dup17_const_fix_32_0_1__0000000000000235_570;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
  wire [31:0] _dup17_const_fix_32_0_1__0000000000000235_801;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
  wire [31:0] _dup17_const_fix_32_0_1__0000000000000235_1032;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
  wire [31:0] _dup17_const_fix_32_0_1__0000000000000235_1263;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
  wire [31:0] _dup17_const_fix_32_0_1__0000000000000235_1494;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
  wire [31:0] _dup17_const_fix_32_0_1__0000000000000235_1725;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
  wire [31:0] _dup17_const_fix_32_0_1__0000000000000235_1956;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
  wire [31:0] _dup17_const_fix_32_0_1__0000000000000235_2320;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
  wire [31:0] _dup17_const_fix_32_0_1__0000000000000235_2684;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
  wire [31:0] _dup17_const_fix_32_0_1__0000000000000235_3048;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
  wire [31:0] _dup17_const_fix_32_0_1__0000000000000235_3412;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
  wire [31:0] _dup17_const_fix_32_0_1__0000000000000235_3776;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
  wire [31:0] _dup17_const_fix_32_0_1__0000000000000235_4140;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
  wire [31:0] _dup17_const_fix_32_0_1__0000000000000235_4504;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
  wire [31:0] _MUL16__dfc_wire_107;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:162:126
  wire [31:0] _dup15_const_fix_32_0_1__0000000000000235_108;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
  wire [31:0] _dup15_const_fix_32_0_1__0000000000000235_339;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
  wire [31:0] _dup15_const_fix_32_0_1__0000000000000235_570;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
  wire [31:0] _dup15_const_fix_32_0_1__0000000000000235_801;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
  wire [31:0] _dup15_const_fix_32_0_1__0000000000000235_1032;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
  wire [31:0] _dup15_const_fix_32_0_1__0000000000000235_1263;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
  wire [31:0] _dup15_const_fix_32_0_1__0000000000000235_1494;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
  wire [31:0] _dup15_const_fix_32_0_1__0000000000000235_1725;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
  wire [31:0] _dup15_const_fix_32_0_1__0000000000000235_1956;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
  wire [31:0] _dup15_const_fix_32_0_1__0000000000000235_2320;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
  wire [31:0] _dup15_const_fix_32_0_1__0000000000000235_2684;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
  wire [31:0] _dup15_const_fix_32_0_1__0000000000000235_3048;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
  wire [31:0] _dup15_const_fix_32_0_1__0000000000000235_3412;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
  wire [31:0] _dup15_const_fix_32_0_1__0000000000000235_3776;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
  wire [31:0] _dup15_const_fix_32_0_1__0000000000000235_4140;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
  wire [31:0] _dup15_const_fix_32_0_1__0000000000000235_4504;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
  wire [31:0] _ADD14__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:160:125
  wire [31:0] _dup13__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:159:106
  wire [31:0] _dup13__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:159:106
  wire [31:0] _dup12__dfc_wire_68_105;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:158:106
  wire [31:0] _dup12__dfc_wire_68_113;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:158:106
  wire [31:0] _ADD11__dfc_wire_100;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:157:125
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_102;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_215;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_227;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_333;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_446;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_458;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_564;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_677;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_689;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_795;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_908;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_920;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_1026;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_1139;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_1151;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_1257;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_1370;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_1382;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_1488;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_1601;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_1613;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_1719;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_1832;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_1844;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_2084;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_2096;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_2448;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_2460;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_2812;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_2824;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_3176;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_3188;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_3540;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_3552;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_3904;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_3916;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_4268;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_4280;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_4632;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _dup10_const_fix_32_0_1__0000000000000080_4644;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
  wire [31:0] _SHL119__dfc_wire_75;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:155:81
  wire [31:0] _CAST8__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:154:76
  wire [31:0] _CAST7__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:153:76
  wire [31:0] _CAST6__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:152:76
  wire [31:0] _CAST5__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:151:76
  wire [31:0] _CAST4__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:150:76
  wire [31:0] _CAST3__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:149:76
  wire [31:0] _CAST2__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:148:76
  wire [31:0] _SHL111__dfc_wire_75;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:147:81
  wire [31:0] _CAST0__dfc_wire_73;	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:146:76

  CAST_1x1_16_32 CAST0 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:146:76
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_4__dfc_wire_45),
    ._dfc_wire_73 (_CAST0__dfc_wire_73)
  );
  SHL11_1x1 SHL111 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:147:81
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_73 (_CAST0__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:146:76
    ._dfc_wire_75 (_SHL111__dfc_wire_75)
  );
  CAST_1x1_16_32 CAST2 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:148:76
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_6__dfc_wire_45),
    ._dfc_wire_73 (_CAST2__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST3 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:149:76
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_2__dfc_wire_45),
    ._dfc_wire_73 (_CAST3__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST4 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:150:76
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_1__dfc_wire_45),
    ._dfc_wire_73 (_CAST4__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST5 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:151:76
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_7__dfc_wire_45),
    ._dfc_wire_73 (_CAST5__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST6 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:152:76
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_5__dfc_wire_45),
    ._dfc_wire_73 (_CAST6__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST7 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:153:76
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_3__dfc_wire_45),
    ._dfc_wire_73 (_CAST7__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST8 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:154:76
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_0__dfc_wire_45),
    ._dfc_wire_73 (_CAST8__dfc_wire_73)
  );
  SHL11_1x1 SHL119 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:155:81
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_73 (_CAST8__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:154:76
    ._dfc_wire_75 (_SHL119__dfc_wire_75)
  );
  dup_1x40 dup10 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .clock                                   (clock),
    .reset                                   (reset),
    .const_fix_32_0_1__0000000000000080      (_const2106_const_fix_32_0_1__0000000000000080),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2163:90
    .const_fix_32_0_1__0000000000000080_102  (_dup10_const_fix_32_0_1__0000000000000080_102),
    .const_fix_32_0_1__0000000000000080_215  (_dup10_const_fix_32_0_1__0000000000000080_215),
    .const_fix_32_0_1__0000000000000080_227  (_dup10_const_fix_32_0_1__0000000000000080_227),
    .const_fix_32_0_1__0000000000000080_333  (_dup10_const_fix_32_0_1__0000000000000080_333),
    .const_fix_32_0_1__0000000000000080_446  (_dup10_const_fix_32_0_1__0000000000000080_446),
    .const_fix_32_0_1__0000000000000080_458  (_dup10_const_fix_32_0_1__0000000000000080_458),
    .const_fix_32_0_1__0000000000000080_564  (_dup10_const_fix_32_0_1__0000000000000080_564),
    .const_fix_32_0_1__0000000000000080_677  (_dup10_const_fix_32_0_1__0000000000000080_677),
    .const_fix_32_0_1__0000000000000080_689  (_dup10_const_fix_32_0_1__0000000000000080_689),
    .const_fix_32_0_1__0000000000000080_795  (_dup10_const_fix_32_0_1__0000000000000080_795),
    .const_fix_32_0_1__0000000000000080_908  (_dup10_const_fix_32_0_1__0000000000000080_908),
    .const_fix_32_0_1__0000000000000080_920  (_dup10_const_fix_32_0_1__0000000000000080_920),
    .const_fix_32_0_1__0000000000000080_1026 (_dup10_const_fix_32_0_1__0000000000000080_1026),
    .const_fix_32_0_1__0000000000000080_1139 (_dup10_const_fix_32_0_1__0000000000000080_1139),
    .const_fix_32_0_1__0000000000000080_1151 (_dup10_const_fix_32_0_1__0000000000000080_1151),
    .const_fix_32_0_1__0000000000000080_1257 (_dup10_const_fix_32_0_1__0000000000000080_1257),
    .const_fix_32_0_1__0000000000000080_1370 (_dup10_const_fix_32_0_1__0000000000000080_1370),
    .const_fix_32_0_1__0000000000000080_1382 (_dup10_const_fix_32_0_1__0000000000000080_1382),
    .const_fix_32_0_1__0000000000000080_1488 (_dup10_const_fix_32_0_1__0000000000000080_1488),
    .const_fix_32_0_1__0000000000000080_1601 (_dup10_const_fix_32_0_1__0000000000000080_1601),
    .const_fix_32_0_1__0000000000000080_1613 (_dup10_const_fix_32_0_1__0000000000000080_1613),
    .const_fix_32_0_1__0000000000000080_1719 (_dup10_const_fix_32_0_1__0000000000000080_1719),
    .const_fix_32_0_1__0000000000000080_1832 (_dup10_const_fix_32_0_1__0000000000000080_1832),
    .const_fix_32_0_1__0000000000000080_1844 (_dup10_const_fix_32_0_1__0000000000000080_1844),
    .const_fix_32_0_1__0000000000000080_2084 (_dup10_const_fix_32_0_1__0000000000000080_2084),
    .const_fix_32_0_1__0000000000000080_2096 (_dup10_const_fix_32_0_1__0000000000000080_2096),
    .const_fix_32_0_1__0000000000000080_2448 (_dup10_const_fix_32_0_1__0000000000000080_2448),
    .const_fix_32_0_1__0000000000000080_2460 (_dup10_const_fix_32_0_1__0000000000000080_2460),
    .const_fix_32_0_1__0000000000000080_2812 (_dup10_const_fix_32_0_1__0000000000000080_2812),
    .const_fix_32_0_1__0000000000000080_2824 (_dup10_const_fix_32_0_1__0000000000000080_2824),
    .const_fix_32_0_1__0000000000000080_3176 (_dup10_const_fix_32_0_1__0000000000000080_3176),
    .const_fix_32_0_1__0000000000000080_3188 (_dup10_const_fix_32_0_1__0000000000000080_3188),
    .const_fix_32_0_1__0000000000000080_3540 (_dup10_const_fix_32_0_1__0000000000000080_3540),
    .const_fix_32_0_1__0000000000000080_3552 (_dup10_const_fix_32_0_1__0000000000000080_3552),
    .const_fix_32_0_1__0000000000000080_3904 (_dup10_const_fix_32_0_1__0000000000000080_3904),
    .const_fix_32_0_1__0000000000000080_3916 (_dup10_const_fix_32_0_1__0000000000000080_3916),
    .const_fix_32_0_1__0000000000000080_4268 (_dup10_const_fix_32_0_1__0000000000000080_4268),
    .const_fix_32_0_1__0000000000000080_4280 (_dup10_const_fix_32_0_1__0000000000000080_4280),
    .const_fix_32_0_1__0000000000000080_4632 (_dup10_const_fix_32_0_1__0000000000000080_4632),
    .const_fix_32_0_1__0000000000000080_4644 (_dup10_const_fix_32_0_1__0000000000000080_4644)
  );
  ADD_2x1 ADD11 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:157:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_SHL119__dfc_wire_75),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:155:81
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_119_3245_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3263:146
    ._dfc_wire_100                          (_ADD11__dfc_wire_100)
  );
  dup_1x2 dup12 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:158:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST4__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:150:76
    ._dfc_wire_68_105 (_dup12__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup12__dfc_wire_68_113)
  );
  dup_1x2 dup13 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:159:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST5__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:151:76
    ._dfc_wire_68_105 (_dup13__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup13__dfc_wire_68_113)
  );
  ADD_2x1 ADD14 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:160:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_12_3244_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3262:142
    .const_fix_32_0_1__0000000000000080_102 (_dup13__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:159:106
    ._dfc_wire_100                          (_ADD14__dfc_wire_100)
  );
  dup_1x16 dup15 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
    .clock                                   (clock),
    .reset                                   (reset),
    .const_fix_32_0_1__0000000000000235      (_const2149_const_fix_32_0_1__0000000000000235),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2167:90
    .const_fix_32_0_1__0000000000000235_108  (_dup15_const_fix_32_0_1__0000000000000235_108),
    .const_fix_32_0_1__0000000000000235_339  (_dup15_const_fix_32_0_1__0000000000000235_339),
    .const_fix_32_0_1__0000000000000235_570  (_dup15_const_fix_32_0_1__0000000000000235_570),
    .const_fix_32_0_1__0000000000000235_801  (_dup15_const_fix_32_0_1__0000000000000235_801),
    .const_fix_32_0_1__0000000000000235_1032 (_dup15_const_fix_32_0_1__0000000000000235_1032),
    .const_fix_32_0_1__0000000000000235_1263 (_dup15_const_fix_32_0_1__0000000000000235_1263),
    .const_fix_32_0_1__0000000000000235_1494 (_dup15_const_fix_32_0_1__0000000000000235_1494),
    .const_fix_32_0_1__0000000000000235_1725 (_dup15_const_fix_32_0_1__0000000000000235_1725),
    .const_fix_32_0_1__0000000000000235_1956 (_dup15_const_fix_32_0_1__0000000000000235_1956),
    .const_fix_32_0_1__0000000000000235_2320 (_dup15_const_fix_32_0_1__0000000000000235_2320),
    .const_fix_32_0_1__0000000000000235_2684 (_dup15_const_fix_32_0_1__0000000000000235_2684),
    .const_fix_32_0_1__0000000000000235_3048 (_dup15_const_fix_32_0_1__0000000000000235_3048),
    .const_fix_32_0_1__0000000000000235_3412 (_dup15_const_fix_32_0_1__0000000000000235_3412),
    .const_fix_32_0_1__0000000000000235_3776 (_dup15_const_fix_32_0_1__0000000000000235_3776),
    .const_fix_32_0_1__0000000000000235_4140 (_dup15_const_fix_32_0_1__0000000000000235_4140),
    .const_fix_32_0_1__0000000000000235_4504 (_dup15_const_fix_32_0_1__0000000000000235_4504)
  );
  MUL_2x1 MUL16 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:162:126
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_70_3243_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3261:142
    ._dfc_wire_104                          (_ADD14__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:160:125
    ._dfc_wire_107                          (_MUL16__dfc_wire_107)
  );
  dup_1x16 dup17 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
    .clock                                   (clock),
    .reset                                   (reset),
    .const_fix_32_0_1__0000000000000235      (_const2074_const_fix_32_0_1__00000000000008e4),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2157:90
    .const_fix_32_0_1__0000000000000235_108  (_dup17_const_fix_32_0_1__0000000000000235_108),
    .const_fix_32_0_1__0000000000000235_339  (_dup17_const_fix_32_0_1__0000000000000235_339),
    .const_fix_32_0_1__0000000000000235_570  (_dup17_const_fix_32_0_1__0000000000000235_570),
    .const_fix_32_0_1__0000000000000235_801  (_dup17_const_fix_32_0_1__0000000000000235_801),
    .const_fix_32_0_1__0000000000000235_1032 (_dup17_const_fix_32_0_1__0000000000000235_1032),
    .const_fix_32_0_1__0000000000000235_1263 (_dup17_const_fix_32_0_1__0000000000000235_1263),
    .const_fix_32_0_1__0000000000000235_1494 (_dup17_const_fix_32_0_1__0000000000000235_1494),
    .const_fix_32_0_1__0000000000000235_1725 (_dup17_const_fix_32_0_1__0000000000000235_1725),
    .const_fix_32_0_1__0000000000000235_1956 (_dup17_const_fix_32_0_1__0000000000000235_1956),
    .const_fix_32_0_1__0000000000000235_2320 (_dup17_const_fix_32_0_1__0000000000000235_2320),
    .const_fix_32_0_1__0000000000000235_2684 (_dup17_const_fix_32_0_1__0000000000000235_2684),
    .const_fix_32_0_1__0000000000000235_3048 (_dup17_const_fix_32_0_1__0000000000000235_3048),
    .const_fix_32_0_1__0000000000000235_3412 (_dup17_const_fix_32_0_1__0000000000000235_3412),
    .const_fix_32_0_1__0000000000000235_3776 (_dup17_const_fix_32_0_1__0000000000000235_3776),
    .const_fix_32_0_1__0000000000000235_4140 (_dup17_const_fix_32_0_1__0000000000000235_4140),
    .const_fix_32_0_1__0000000000000235_4504 (_dup17_const_fix_32_0_1__0000000000000235_4504)
  );
  MUL_2x1 MUL18 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:164:126
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_34_3242_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3260:142
    ._dfc_wire_104                          (_dup12__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:158:106
    ._dfc_wire_107                          (_MUL18__dfc_wire_107)
  );
  dup_1x2 dup19 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:165:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL16__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:162:126
    ._dfc_wire_68_105 (_dup19__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup19__dfc_wire_68_113)
  );
  ADD_2x1 ADD20 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:166:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup19__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:165:106
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_167_3241_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3259:146
    ._dfc_wire_100                          (_ADD20__dfc_wire_100)
  );
  dup_1x16 dup21 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
    .clock                                   (clock),
    .reset                                   (reset),
    .const_fix_32_0_1__0000000000000235      (_const2081_const_fix_32_0_1__0000000000000d4e),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2158:90
    .const_fix_32_0_1__0000000000000235_108  (_dup21_const_fix_32_0_1__0000000000000235_108),
    .const_fix_32_0_1__0000000000000235_339  (_dup21_const_fix_32_0_1__0000000000000235_339),
    .const_fix_32_0_1__0000000000000235_570  (_dup21_const_fix_32_0_1__0000000000000235_570),
    .const_fix_32_0_1__0000000000000235_801  (_dup21_const_fix_32_0_1__0000000000000235_801),
    .const_fix_32_0_1__0000000000000235_1032 (_dup21_const_fix_32_0_1__0000000000000235_1032),
    .const_fix_32_0_1__0000000000000235_1263 (_dup21_const_fix_32_0_1__0000000000000235_1263),
    .const_fix_32_0_1__0000000000000235_1494 (_dup21_const_fix_32_0_1__0000000000000235_1494),
    .const_fix_32_0_1__0000000000000235_1725 (_dup21_const_fix_32_0_1__0000000000000235_1725),
    .const_fix_32_0_1__0000000000000235_1956 (_dup21_const_fix_32_0_1__0000000000000235_1956),
    .const_fix_32_0_1__0000000000000235_2320 (_dup21_const_fix_32_0_1__0000000000000235_2320),
    .const_fix_32_0_1__0000000000000235_2684 (_dup21_const_fix_32_0_1__0000000000000235_2684),
    .const_fix_32_0_1__0000000000000235_3048 (_dup21_const_fix_32_0_1__0000000000000235_3048),
    .const_fix_32_0_1__0000000000000235_3412 (_dup21_const_fix_32_0_1__0000000000000235_3412),
    .const_fix_32_0_1__0000000000000235_3776 (_dup21_const_fix_32_0_1__0000000000000235_3776),
    .const_fix_32_0_1__0000000000000235_4140 (_dup21_const_fix_32_0_1__0000000000000235_4140),
    .const_fix_32_0_1__0000000000000235_4504 (_dup21_const_fix_32_0_1__0000000000000235_4504)
  );
  MUL_2x1 MUL22 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:168:126
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_90_3238_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3256:142
    ._dfc_wire_104                          (_dup13__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:159:106
    ._dfc_wire_107                          (_MUL22__dfc_wire_107)
  );
  SUB_2x1 SUB23 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:169:104
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup19__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:165:106
    ._dfc_wire_118    (_delay_fixed_32_0_1_93_3236_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3254:142
    ._dfc_wire_121    (_SUB23__dfc_wire_121)
  );
  dup_1x2 dup24 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:170:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST6__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:152:76
    ._dfc_wire_68_105 (_dup24__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup24__dfc_wire_68_113)
  );
  dup_1x2 dup25 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:171:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST7__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:153:76
    ._dfc_wire_68_105 (_dup25__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup25__dfc_wire_68_113)
  );
  ADD_2x1 ADD26 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:172:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup24__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:170:106
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_140_3233_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3251:146
    ._dfc_wire_100                          (_ADD26__dfc_wire_100)
  );
  dup_1x16 dup27 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
    .clock                                   (clock),
    .reset                                   (reset),
    .const_fix_32_0_1__0000000000000235      (_const2097_const_fix_32_0_1__0000000000000968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2160:90
    .const_fix_32_0_1__0000000000000235_108  (_dup27_const_fix_32_0_1__0000000000000235_108),
    .const_fix_32_0_1__0000000000000235_339  (_dup27_const_fix_32_0_1__0000000000000235_339),
    .const_fix_32_0_1__0000000000000235_570  (_dup27_const_fix_32_0_1__0000000000000235_570),
    .const_fix_32_0_1__0000000000000235_801  (_dup27_const_fix_32_0_1__0000000000000235_801),
    .const_fix_32_0_1__0000000000000235_1032 (_dup27_const_fix_32_0_1__0000000000000235_1032),
    .const_fix_32_0_1__0000000000000235_1263 (_dup27_const_fix_32_0_1__0000000000000235_1263),
    .const_fix_32_0_1__0000000000000235_1494 (_dup27_const_fix_32_0_1__0000000000000235_1494),
    .const_fix_32_0_1__0000000000000235_1725 (_dup27_const_fix_32_0_1__0000000000000235_1725),
    .const_fix_32_0_1__0000000000000235_1956 (_dup27_const_fix_32_0_1__0000000000000235_1956),
    .const_fix_32_0_1__0000000000000235_2320 (_dup27_const_fix_32_0_1__0000000000000235_2320),
    .const_fix_32_0_1__0000000000000235_2684 (_dup27_const_fix_32_0_1__0000000000000235_2684),
    .const_fix_32_0_1__0000000000000235_3048 (_dup27_const_fix_32_0_1__0000000000000235_3048),
    .const_fix_32_0_1__0000000000000235_3412 (_dup27_const_fix_32_0_1__0000000000000235_3412),
    .const_fix_32_0_1__0000000000000235_3776 (_dup27_const_fix_32_0_1__0000000000000235_3776),
    .const_fix_32_0_1__0000000000000235_4140 (_dup27_const_fix_32_0_1__0000000000000235_4140),
    .const_fix_32_0_1__0000000000000235_4504 (_dup27_const_fix_32_0_1__0000000000000235_4504)
  );
  MUL_2x1 MUL28 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:174:126
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_230_3231_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3249:146
    ._dfc_wire_104                          (_ADD26__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:172:125
    ._dfc_wire_107                          (_MUL28__dfc_wire_107)
  );
  dup_1x16 dup29 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
    .clock                                   (clock),
    .reset                                   (reset),
    .const_fix_32_0_1__0000000000000235      (_const2065_const_fix_32_0_1__000000000000031f),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2155:90
    .const_fix_32_0_1__0000000000000235_108  (_dup29_const_fix_32_0_1__0000000000000235_108),
    .const_fix_32_0_1__0000000000000235_339  (_dup29_const_fix_32_0_1__0000000000000235_339),
    .const_fix_32_0_1__0000000000000235_570  (_dup29_const_fix_32_0_1__0000000000000235_570),
    .const_fix_32_0_1__0000000000000235_801  (_dup29_const_fix_32_0_1__0000000000000235_801),
    .const_fix_32_0_1__0000000000000235_1032 (_dup29_const_fix_32_0_1__0000000000000235_1032),
    .const_fix_32_0_1__0000000000000235_1263 (_dup29_const_fix_32_0_1__0000000000000235_1263),
    .const_fix_32_0_1__0000000000000235_1494 (_dup29_const_fix_32_0_1__0000000000000235_1494),
    .const_fix_32_0_1__0000000000000235_1725 (_dup29_const_fix_32_0_1__0000000000000235_1725),
    .const_fix_32_0_1__0000000000000235_1956 (_dup29_const_fix_32_0_1__0000000000000235_1956),
    .const_fix_32_0_1__0000000000000235_2320 (_dup29_const_fix_32_0_1__0000000000000235_2320),
    .const_fix_32_0_1__0000000000000235_2684 (_dup29_const_fix_32_0_1__0000000000000235_2684),
    .const_fix_32_0_1__0000000000000235_3048 (_dup29_const_fix_32_0_1__0000000000000235_3048),
    .const_fix_32_0_1__0000000000000235_3412 (_dup29_const_fix_32_0_1__0000000000000235_3412),
    .const_fix_32_0_1__0000000000000235_3776 (_dup29_const_fix_32_0_1__0000000000000235_3776),
    .const_fix_32_0_1__0000000000000235_4140 (_dup29_const_fix_32_0_1__0000000000000235_4140),
    .const_fix_32_0_1__0000000000000235_4504 (_dup29_const_fix_32_0_1__0000000000000235_4504)
  );
  MUL_2x1 MUL30 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:176:126
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_72_3227_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3245:142
    ._dfc_wire_104                          (_dup24__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:170:106
    ._dfc_wire_107                          (_MUL30__dfc_wire_107)
  );
  dup_1x2 dup31 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:177:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL28__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:174:126
    ._dfc_wire_68_105 (_dup31__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup31__dfc_wire_68_113)
  );
  SUB_2x1 SUB32 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:178:104
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup31__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:177:106
    ._dfc_wire_118    (_delay_fixed_32_0_1_148_3226_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3244:146
    ._dfc_wire_121    (_SUB32__dfc_wire_121)
  );
  dup_1x16 dup33 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
    .clock                                   (clock),
    .reset                                   (reset),
    .const_fix_32_0_1__0000000000000235      (_const2068_const_fix_32_0_1__0000000000000fb1),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2156:90
    .const_fix_32_0_1__0000000000000235_108  (_dup33_const_fix_32_0_1__0000000000000235_108),
    .const_fix_32_0_1__0000000000000235_339  (_dup33_const_fix_32_0_1__0000000000000235_339),
    .const_fix_32_0_1__0000000000000235_570  (_dup33_const_fix_32_0_1__0000000000000235_570),
    .const_fix_32_0_1__0000000000000235_801  (_dup33_const_fix_32_0_1__0000000000000235_801),
    .const_fix_32_0_1__0000000000000235_1032 (_dup33_const_fix_32_0_1__0000000000000235_1032),
    .const_fix_32_0_1__0000000000000235_1263 (_dup33_const_fix_32_0_1__0000000000000235_1263),
    .const_fix_32_0_1__0000000000000235_1494 (_dup33_const_fix_32_0_1__0000000000000235_1494),
    .const_fix_32_0_1__0000000000000235_1725 (_dup33_const_fix_32_0_1__0000000000000235_1725),
    .const_fix_32_0_1__0000000000000235_1956 (_dup33_const_fix_32_0_1__0000000000000235_1956),
    .const_fix_32_0_1__0000000000000235_2320 (_dup33_const_fix_32_0_1__0000000000000235_2320),
    .const_fix_32_0_1__0000000000000235_2684 (_dup33_const_fix_32_0_1__0000000000000235_2684),
    .const_fix_32_0_1__0000000000000235_3048 (_dup33_const_fix_32_0_1__0000000000000235_3048),
    .const_fix_32_0_1__0000000000000235_3412 (_dup33_const_fix_32_0_1__0000000000000235_3412),
    .const_fix_32_0_1__0000000000000235_3776 (_dup33_const_fix_32_0_1__0000000000000235_3776),
    .const_fix_32_0_1__0000000000000235_4140 (_dup33_const_fix_32_0_1__0000000000000235_4140),
    .const_fix_32_0_1__0000000000000235_4504 (_dup33_const_fix_32_0_1__0000000000000235_4504)
  );
  MUL_2x1 MUL34 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:180:126
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_dup33_const_fix_32_0_1__0000000000000235_108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
    ._dfc_wire_104                          (_delay_fixed_32_0_1_10_3224_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3242:142
    ._dfc_wire_107                          (_MUL34__dfc_wire_107)
  );
  SUB_2x1 SUB35 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:181:104
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup31__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:177:106
    ._dfc_wire_118    (_delay_fixed_32_0_1_280_3223_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3241:146
    ._dfc_wire_121    (_SUB35__dfc_wire_121)
  );
  dup_1x2 dup36 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:182:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD11__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:157:125
    ._dfc_wire_68_105 (_dup36__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup36__dfc_wire_68_113)
  );
  dup_1x2 dup37 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:183:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHL111__dfc_wire_75),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:147:81
    ._dfc_wire_68_105 (_dup37__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup37__dfc_wire_68_113)
  );
  ADD_2x1 ADD38 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:184:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup36__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:182:106
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_5_3219_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3237:138
    ._dfc_wire_100                          (_ADD38__dfc_wire_100)
  );
  SUB_2x1 SUB39 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:185:104
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup36__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:182:106
    ._dfc_wire_118    (_delay_fixed_32_0_1_5_3217_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3235:138
    ._dfc_wire_121    (_SUB39__dfc_wire_121)
  );
  dup_1x2 dup40 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:186:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST3__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:149:76
    ._dfc_wire_68_105 (_dup40__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup40__dfc_wire_68_113)
  );
  dup_1x2 dup41 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:187:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST2__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:148:76
    ._dfc_wire_68_105 (_dup41__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup41__dfc_wire_68_113)
  );
  ADD_2x1 ADD42 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:188:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup40__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:186:106
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1_3213_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3231:138
    ._dfc_wire_100                          (_ADD42__dfc_wire_100)
  );
  dup_1x16 dup43 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
    .clock                                   (clock),
    .reset                                   (reset),
    .const_fix_32_0_1__0000000000000235      (_const2111_const_fix_32_0_1__0000000000000454),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2164:90
    .const_fix_32_0_1__0000000000000235_108  (_dup43_const_fix_32_0_1__0000000000000235_108),
    .const_fix_32_0_1__0000000000000235_339  (_dup43_const_fix_32_0_1__0000000000000235_339),
    .const_fix_32_0_1__0000000000000235_570  (_dup43_const_fix_32_0_1__0000000000000235_570),
    .const_fix_32_0_1__0000000000000235_801  (_dup43_const_fix_32_0_1__0000000000000235_801),
    .const_fix_32_0_1__0000000000000235_1032 (_dup43_const_fix_32_0_1__0000000000000235_1032),
    .const_fix_32_0_1__0000000000000235_1263 (_dup43_const_fix_32_0_1__0000000000000235_1263),
    .const_fix_32_0_1__0000000000000235_1494 (_dup43_const_fix_32_0_1__0000000000000235_1494),
    .const_fix_32_0_1__0000000000000235_1725 (_dup43_const_fix_32_0_1__0000000000000235_1725),
    .const_fix_32_0_1__0000000000000235_1956 (_dup43_const_fix_32_0_1__0000000000000235_1956),
    .const_fix_32_0_1__0000000000000235_2320 (_dup43_const_fix_32_0_1__0000000000000235_2320),
    .const_fix_32_0_1__0000000000000235_2684 (_dup43_const_fix_32_0_1__0000000000000235_2684),
    .const_fix_32_0_1__0000000000000235_3048 (_dup43_const_fix_32_0_1__0000000000000235_3048),
    .const_fix_32_0_1__0000000000000235_3412 (_dup43_const_fix_32_0_1__0000000000000235_3412),
    .const_fix_32_0_1__0000000000000235_3776 (_dup43_const_fix_32_0_1__0000000000000235_3776),
    .const_fix_32_0_1__0000000000000235_4140 (_dup43_const_fix_32_0_1__0000000000000235_4140),
    .const_fix_32_0_1__0000000000000235_4504 (_dup43_const_fix_32_0_1__0000000000000235_4504)
  );
  MUL_2x1 MUL44 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:190:126
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_188_3209_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3227:146
    ._dfc_wire_104                          (_ADD42__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:188:125
    ._dfc_wire_107                          (_MUL44__dfc_wire_107)
  );
  dup_1x16 dup45 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
    .clock                                   (clock),
    .reset                                   (reset),
    .const_fix_32_0_1__0000000000000235      (_const2098_const_fix_32_0_1__0000000000000ec8),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2161:90
    .const_fix_32_0_1__0000000000000235_108  (_dup45_const_fix_32_0_1__0000000000000235_108),
    .const_fix_32_0_1__0000000000000235_339  (_dup45_const_fix_32_0_1__0000000000000235_339),
    .const_fix_32_0_1__0000000000000235_570  (_dup45_const_fix_32_0_1__0000000000000235_570),
    .const_fix_32_0_1__0000000000000235_801  (_dup45_const_fix_32_0_1__0000000000000235_801),
    .const_fix_32_0_1__0000000000000235_1032 (_dup45_const_fix_32_0_1__0000000000000235_1032),
    .const_fix_32_0_1__0000000000000235_1263 (_dup45_const_fix_32_0_1__0000000000000235_1263),
    .const_fix_32_0_1__0000000000000235_1494 (_dup45_const_fix_32_0_1__0000000000000235_1494),
    .const_fix_32_0_1__0000000000000235_1725 (_dup45_const_fix_32_0_1__0000000000000235_1725),
    .const_fix_32_0_1__0000000000000235_1956 (_dup45_const_fix_32_0_1__0000000000000235_1956),
    .const_fix_32_0_1__0000000000000235_2320 (_dup45_const_fix_32_0_1__0000000000000235_2320),
    .const_fix_32_0_1__0000000000000235_2684 (_dup45_const_fix_32_0_1__0000000000000235_2684),
    .const_fix_32_0_1__0000000000000235_3048 (_dup45_const_fix_32_0_1__0000000000000235_3048),
    .const_fix_32_0_1__0000000000000235_3412 (_dup45_const_fix_32_0_1__0000000000000235_3412),
    .const_fix_32_0_1__0000000000000235_3776 (_dup45_const_fix_32_0_1__0000000000000235_3776),
    .const_fix_32_0_1__0000000000000235_4140 (_dup45_const_fix_32_0_1__0000000000000235_4140),
    .const_fix_32_0_1__0000000000000235_4504 (_dup45_const_fix_32_0_1__0000000000000235_4504)
  );
  MUL_2x1 MUL46 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:192:126
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_100_3208_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3226:146
    ._dfc_wire_104                          (_dup41__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:187:106
    ._dfc_wire_107                          (_MUL46__dfc_wire_107)
  );
  dup_1x2 dup47 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:193:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL44__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:190:126
    ._dfc_wire_68_105 (_dup47__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup47__dfc_wire_68_113)
  );
  SUB_2x1 SUB48 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:194:104
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup47__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:193:106
    ._dfc_wire_118    (_delay_fixed_32_0_1_85_3207_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3225:142
    ._dfc_wire_121    (_SUB48__dfc_wire_121)
  );
  dup_1x16 dup49 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
    .clock                                   (clock),
    .reset                                   (reset),
    .const_fix_32_0_1__0000000000000235      (_const2060_const_fix_32_0_1__0000000000000620),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2154:90
    .const_fix_32_0_1__0000000000000235_108  (_dup49_const_fix_32_0_1__0000000000000235_108),
    .const_fix_32_0_1__0000000000000235_339  (_dup49_const_fix_32_0_1__0000000000000235_339),
    .const_fix_32_0_1__0000000000000235_570  (_dup49_const_fix_32_0_1__0000000000000235_570),
    .const_fix_32_0_1__0000000000000235_801  (_dup49_const_fix_32_0_1__0000000000000235_801),
    .const_fix_32_0_1__0000000000000235_1032 (_dup49_const_fix_32_0_1__0000000000000235_1032),
    .const_fix_32_0_1__0000000000000235_1263 (_dup49_const_fix_32_0_1__0000000000000235_1263),
    .const_fix_32_0_1__0000000000000235_1494 (_dup49_const_fix_32_0_1__0000000000000235_1494),
    .const_fix_32_0_1__0000000000000235_1725 (_dup49_const_fix_32_0_1__0000000000000235_1725),
    .const_fix_32_0_1__0000000000000235_1956 (_dup49_const_fix_32_0_1__0000000000000235_1956),
    .const_fix_32_0_1__0000000000000235_2320 (_dup49_const_fix_32_0_1__0000000000000235_2320),
    .const_fix_32_0_1__0000000000000235_2684 (_dup49_const_fix_32_0_1__0000000000000235_2684),
    .const_fix_32_0_1__0000000000000235_3048 (_dup49_const_fix_32_0_1__0000000000000235_3048),
    .const_fix_32_0_1__0000000000000235_3412 (_dup49_const_fix_32_0_1__0000000000000235_3412),
    .const_fix_32_0_1__0000000000000235_3776 (_dup49_const_fix_32_0_1__0000000000000235_3776),
    .const_fix_32_0_1__0000000000000235_4140 (_dup49_const_fix_32_0_1__0000000000000235_4140),
    .const_fix_32_0_1__0000000000000235_4504 (_dup49_const_fix_32_0_1__0000000000000235_4504)
  );
  MUL_2x1 MUL50 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:196:126
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_157_3205_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3223:146
    ._dfc_wire_104                          (_dup40__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:186:106
    ._dfc_wire_107                          (_MUL50__dfc_wire_107)
  );
  ADD_2x1 ADD51 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:197:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup47__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:193:106
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_77_3204_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3222:142
    ._dfc_wire_100                          (_ADD51__dfc_wire_100)
  );
  dup_1x2 dup52 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:198:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD20__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:166:125
    ._dfc_wire_68_105 (_dup52__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup52__dfc_wire_68_113)
  );
  dup_1x2 dup53 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:199:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB32__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:178:104
    ._dfc_wire_68_105 (_dup53__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup53__dfc_wire_68_113)
  );
  ADD_2x1 ADD54 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:200:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_11_3201_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3219:142
    .const_fix_32_0_1__0000000000000080_102 (_dup53__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:199:106
    ._dfc_wire_100                          (_ADD54__dfc_wire_100)
  );
  SUB_2x1 SUB55 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:201:104
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_11_3200_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3218:142
    ._dfc_wire_118    (_dup53__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:199:106
    ._dfc_wire_121    (_SUB55__dfc_wire_121)
  );
  dup_1x2 dup56 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:202:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB23__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:169:104
    ._dfc_wire_68_105 (_dup56__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup56__dfc_wire_68_113)
  );
  dup_1x2 dup57 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:203:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB35__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:181:104
    ._dfc_wire_68_105 (_dup57__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup57__dfc_wire_68_113)
  );
  ADD_2x1 ADD58 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:204:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_22_3195_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3213:142
    .const_fix_32_0_1__0000000000000080_102 (_dup57__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:203:106
    ._dfc_wire_100                          (_ADD58__dfc_wire_100)
  );
  SUB_2x1 SUB59 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:205:104
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_22_3192_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3210:142
    ._dfc_wire_118    (_dup57__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:203:106
    ._dfc_wire_121    (_SUB59__dfc_wire_121)
  );
  dup_1x2 dup60 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:206:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD38__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:184:125
    ._dfc_wire_68_105 (_dup60__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup60__dfc_wire_68_113)
  );
  dup_1x2 dup61 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:207:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD51__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:197:125
    ._dfc_wire_68_105 (_dup61__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup61__dfc_wire_68_113)
  );
  ADD_2x1 ADD62 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:208:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_178_3191_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3209:146
    .const_fix_32_0_1__0000000000000080_102 (_dup61__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:207:106
    ._dfc_wire_100                          (_ADD62__dfc_wire_100)
  );
  SUB_2x1 SUB63 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:209:104
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_178_3190_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3208:146
    ._dfc_wire_118    (_dup61__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:207:106
    ._dfc_wire_121    (_SUB63__dfc_wire_121)
  );
  dup_1x2 dup64 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:210:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB39__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:185:104
    ._dfc_wire_68_105 (_dup64__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup64__dfc_wire_68_113)
  );
  dup_1x2 dup65 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:211:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB48__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:194:104
    ._dfc_wire_68_105 (_dup65__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup65__dfc_wire_68_113)
  );
  ADD_2x1 ADD66 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:212:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_205_3189_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3207:146
    .const_fix_32_0_1__0000000000000080_102 (_dup65__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:211:106
    ._dfc_wire_100                          (_ADD66__dfc_wire_100)
  );
  SUB_2x1 SUB67 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:213:104
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_205_3188_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3206:146
    ._dfc_wire_118    (_dup65__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:211:106
    ._dfc_wire_121    (_SUB67__dfc_wire_121)
  );
  dup_1x2 dup68 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:214:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB55__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:201:104
    ._dfc_wire_68_105 (_dup68__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup68__dfc_wire_68_113)
  );
  dup_1x2 dup69 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:215:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB59__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:205:104
    ._dfc_wire_68_105 (_dup69__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup69__dfc_wire_68_113)
  );
  ADD_2x1 ADD70 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:216:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup68__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:214:106
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1_3187_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3205:138
    ._dfc_wire_100                          (_ADD70__dfc_wire_100)
  );
  dup_1x32 dup71 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .clock                                   (clock),
    .reset                                   (reset),
    .const_fix_32_0_1__00000000000000b5      (_const2102_const_fix_32_0_1__00000000000000b5),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2162:90
    .const_fix_32_0_1__00000000000000b5_211  (_dup71_const_fix_32_0_1__00000000000000b5_211),
    .const_fix_32_0_1__00000000000000b5_223  (_dup71_const_fix_32_0_1__00000000000000b5_223),
    .const_fix_32_0_1__00000000000000b5_442  (_dup71_const_fix_32_0_1__00000000000000b5_442),
    .const_fix_32_0_1__00000000000000b5_454  (_dup71_const_fix_32_0_1__00000000000000b5_454),
    .const_fix_32_0_1__00000000000000b5_673  (_dup71_const_fix_32_0_1__00000000000000b5_673),
    .const_fix_32_0_1__00000000000000b5_685  (_dup71_const_fix_32_0_1__00000000000000b5_685),
    .const_fix_32_0_1__00000000000000b5_904  (_dup71_const_fix_32_0_1__00000000000000b5_904),
    .const_fix_32_0_1__00000000000000b5_916  (_dup71_const_fix_32_0_1__00000000000000b5_916),
    .const_fix_32_0_1__00000000000000b5_1135 (_dup71_const_fix_32_0_1__00000000000000b5_1135),
    .const_fix_32_0_1__00000000000000b5_1147 (_dup71_const_fix_32_0_1__00000000000000b5_1147),
    .const_fix_32_0_1__00000000000000b5_1366 (_dup71_const_fix_32_0_1__00000000000000b5_1366),
    .const_fix_32_0_1__00000000000000b5_1378 (_dup71_const_fix_32_0_1__00000000000000b5_1378),
    .const_fix_32_0_1__00000000000000b5_1597 (_dup71_const_fix_32_0_1__00000000000000b5_1597),
    .const_fix_32_0_1__00000000000000b5_1609 (_dup71_const_fix_32_0_1__00000000000000b5_1609),
    .const_fix_32_0_1__00000000000000b5_1828 (_dup71_const_fix_32_0_1__00000000000000b5_1828),
    .const_fix_32_0_1__00000000000000b5_1840 (_dup71_const_fix_32_0_1__00000000000000b5_1840),
    .const_fix_32_0_1__00000000000000b5_2080 (_dup71_const_fix_32_0_1__00000000000000b5_2080),
    .const_fix_32_0_1__00000000000000b5_2092 (_dup71_const_fix_32_0_1__00000000000000b5_2092),
    .const_fix_32_0_1__00000000000000b5_2444 (_dup71_const_fix_32_0_1__00000000000000b5_2444),
    .const_fix_32_0_1__00000000000000b5_2456 (_dup71_const_fix_32_0_1__00000000000000b5_2456),
    .const_fix_32_0_1__00000000000000b5_2808 (_dup71_const_fix_32_0_1__00000000000000b5_2808),
    .const_fix_32_0_1__00000000000000b5_2820 (_dup71_const_fix_32_0_1__00000000000000b5_2820),
    .const_fix_32_0_1__00000000000000b5_3172 (_dup71_const_fix_32_0_1__00000000000000b5_3172),
    .const_fix_32_0_1__00000000000000b5_3184 (_dup71_const_fix_32_0_1__00000000000000b5_3184),
    .const_fix_32_0_1__00000000000000b5_3536 (_dup71_const_fix_32_0_1__00000000000000b5_3536),
    .const_fix_32_0_1__00000000000000b5_3548 (_dup71_const_fix_32_0_1__00000000000000b5_3548),
    .const_fix_32_0_1__00000000000000b5_3900 (_dup71_const_fix_32_0_1__00000000000000b5_3900),
    .const_fix_32_0_1__00000000000000b5_3912 (_dup71_const_fix_32_0_1__00000000000000b5_3912),
    .const_fix_32_0_1__00000000000000b5_4264 (_dup71_const_fix_32_0_1__00000000000000b5_4264),
    .const_fix_32_0_1__00000000000000b5_4276 (_dup71_const_fix_32_0_1__00000000000000b5_4276),
    .const_fix_32_0_1__00000000000000b5_4628 (_dup71_const_fix_32_0_1__00000000000000b5_4628),
    .const_fix_32_0_1__00000000000000b5_4640 (_dup71_const_fix_32_0_1__00000000000000b5_4640)
  );
  MUL_2x1 MUL72 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:218:126
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_484_3186_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3204:146
    ._dfc_wire_104                          (_ADD70__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:216:125
    ._dfc_wire_107                          (_MUL72__dfc_wire_107)
  );
  ADD_2x1 ADD73 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:219:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL72__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:218:126
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_566_3185_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3203:146
    ._dfc_wire_100                          (_ADD73__dfc_wire_100)
  );
  SHR8_1x1 SHR874 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:220:83
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD73__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:219:125
    ._dfc_wire_216 (_SHR874__dfc_wire_216)
  );
  SUB_2x1 SUB75 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:221:104
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup68__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:214:106
    ._dfc_wire_118    (_delay_fixed_32_0_1_1_3184_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3202:138
    ._dfc_wire_121    (_SUB75__dfc_wire_121)
  );
  MUL_2x1 MUL76 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:222:126
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_461_3183_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3201:146
    ._dfc_wire_104                          (_SUB75__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:221:104
    ._dfc_wire_107                          (_MUL76__dfc_wire_107)
  );
  ADD_2x1 ADD77 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:223:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL76__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:222:126
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_552_3182_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3200:146
    ._dfc_wire_100                          (_ADD77__dfc_wire_100)
  );
  SHR8_1x1 SHR878 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:224:83
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD77__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:223:125
    ._dfc_wire_216 (_SHR878__dfc_wire_216)
  );
  dup_1x2 dup79 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:225:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD62__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:208:125
    ._dfc_wire_68_105 (_dup79__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup79__dfc_wire_68_113)
  );
  dup_1x2 dup80 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:226:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD54__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:200:125
    ._dfc_wire_68_105 (_dup80__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup80__dfc_wire_68_113)
  );
  ADD_2x1 ADD81 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:227:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_46_3181_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3199:142
    .const_fix_32_0_1__0000000000000080_102 (_dup80__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:226:106
    ._dfc_wire_100                          (_ADD81__dfc_wire_100)
  );
  SHR8_1x1 SHR882 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:228:83
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD81__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:227:125
    ._dfc_wire_216 (_SHR882__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST83 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:229:83
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR882__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:228:83
    ._dfc_wire_236 (_CAST83__dfc_wire_236)
  );
  dup_1x2 dup84 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:230:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD66__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:212:125
    ._dfc_wire_68_105 (_dup84__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup84__dfc_wire_68_113)
  );
  dup_1x2 dup85 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:231:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR874__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:220:83
    ._dfc_wire_68_105 (_dup85__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup85__dfc_wire_68_113)
  );
  ADD_2x1 ADD86 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:232:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_232_3180_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3198:146
    .const_fix_32_0_1__0000000000000080_102 (_dup85__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:231:106
    ._dfc_wire_100                          (_ADD86__dfc_wire_100)
  );
  SHR8_1x1 SHR887 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:233:83
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD86__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:232:125
    ._dfc_wire_216 (_SHR887__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST88 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:234:83
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR887__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:233:83
    ._dfc_wire_236 (_CAST88__dfc_wire_236)
  );
  dup_1x2 dup89 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:235:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB67__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:213:104
    ._dfc_wire_68_105 (_dup89__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup89__dfc_wire_68_113)
  );
  dup_1x2 dup90 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:236:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR878__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:224:83
    ._dfc_wire_68_105 (_dup90__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup90__dfc_wire_68_113)
  );
  ADD_2x1 ADD91 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:237:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_139_3179_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3197:146
    .const_fix_32_0_1__0000000000000080_102 (_dup90__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:236:106
    ._dfc_wire_100                          (_ADD91__dfc_wire_100)
  );
  SHR8_1x1 SHR892 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:238:83
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD91__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:237:125
    ._dfc_wire_216 (_SHR892__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST93 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:239:83
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR892__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:238:83
    ._dfc_wire_236 (_CAST93__dfc_wire_236)
  );
  dup_1x2 dup94 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:240:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB63__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:209:104
    ._dfc_wire_68_105 (_dup94__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup94__dfc_wire_68_113)
  );
  dup_1x2 dup95 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:241:106
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD58__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:204:125
    ._dfc_wire_68_105 (_dup95__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup95__dfc_wire_68_113)
  );
  ADD_2x1 ADD96 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:242:125
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_81_3178_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3196:142
    .const_fix_32_0_1__0000000000000080_102 (_dup95__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:241:106
    ._dfc_wire_100                          (_ADD96__dfc_wire_100)
  );
  SHR8_1x1 SHR897 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:243:83
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD96__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:242:125
    ._dfc_wire_216 (_SHR897__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST98 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:244:83
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR897__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:243:83
    ._dfc_wire_236 (_CAST98__dfc_wire_236)
  );
  SUB_2x1 SUB99 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:245:104
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_81_3177_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3195:142
    ._dfc_wire_118    (_dup95__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:241:106
    ._dfc_wire_121    (_SUB99__dfc_wire_121)
  );
  SHR8_1x1 SHR8100 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:246:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB99__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:245:104
    ._dfc_wire_216 (_SHR8100__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST101 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:247:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8100__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:246:87
    ._dfc_wire_236 (_CAST101__dfc_wire_236)
  );
  SUB_2x1 SUB102 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:248:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_139_3174_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3192:146
    ._dfc_wire_118    (_dup90__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:236:106
    ._dfc_wire_121    (_SUB102__dfc_wire_121)
  );
  SHR8_1x1 SHR8103 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:249:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB102__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:248:109
    ._dfc_wire_216 (_SHR8103__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST104 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:250:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8103__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:249:87
    ._dfc_wire_236 (_CAST104__dfc_wire_236)
  );
  SUB_2x1 SUB105 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:251:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_232_3172_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3190:146
    ._dfc_wire_118    (_dup85__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:231:106
    ._dfc_wire_121    (_SUB105__dfc_wire_121)
  );
  SHR8_1x1 SHR8106 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:252:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB105__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:251:109
    ._dfc_wire_216 (_SHR8106__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST107 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:253:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8106__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:252:87
    ._dfc_wire_236 (_CAST107__dfc_wire_236)
  );
  SUB_2x1 SUB108 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:254:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_46_3170_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3188:142
    ._dfc_wire_118    (_dup80__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:226:106
    ._dfc_wire_121    (_SUB108__dfc_wire_121)
  );
  SHR8_1x1 SHR8109 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:255:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB108__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:254:109
    ._dfc_wire_216 (_SHR8109__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST110 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:256:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8109__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:255:87
    ._dfc_wire_236 (_CAST110__dfc_wire_236)
  );
  CAST_1x1_16_32 CAST111 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:257:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_12__dfc_wire_45),
    ._dfc_wire_73 (_CAST111__dfc_wire_73)
  );
  SHL11_1x1 SHL11112 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:258:89
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_73 (_CAST111__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:257:84
    ._dfc_wire_75 (_SHL11112__dfc_wire_75)
  );
  CAST_1x1_16_32 CAST113 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:259:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_14__dfc_wire_45),
    ._dfc_wire_73 (_CAST113__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST114 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:260:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_10__dfc_wire_45),
    ._dfc_wire_73 (_CAST114__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST115 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:261:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_9__dfc_wire_45),
    ._dfc_wire_73 (_CAST115__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST116 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:262:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_15__dfc_wire_45),
    ._dfc_wire_73 (_CAST116__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST117 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:263:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_13__dfc_wire_45),
    ._dfc_wire_73 (_CAST117__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST118 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:264:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_11__dfc_wire_45),
    ._dfc_wire_73 (_CAST118__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST119 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:265:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_8__dfc_wire_45),
    ._dfc_wire_73 (_CAST119__dfc_wire_73)
  );
  SHL11_1x1 SHL11120 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:266:89
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_73 (_CAST119__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:265:84
    ._dfc_wire_75 (_SHL11120__dfc_wire_75)
  );
  ADD_2x1 ADD121 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:267:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_SHL11120__dfc_wire_75),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:266:89
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_113_3157_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3175:146
    ._dfc_wire_100                          (_ADD121__dfc_wire_100)
  );
  dup_1x2 dup122 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:268:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST115__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:261:84
    ._dfc_wire_68_105 (_dup122__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup122__dfc_wire_68_113)
  );
  dup_1x2 dup123 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:269:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST116__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:262:84
    ._dfc_wire_68_105 (_dup123__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup123__dfc_wire_68_113)
  );
  ADD_2x1 ADD124 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:270:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_54_3155_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3173:142
    .const_fix_32_0_1__0000000000000080_102 (_dup123__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:269:111
    ._dfc_wire_100                          (_ADD124__dfc_wire_100)
  );
  MUL_2x1 MUL125 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:271:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_73_3154_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3172:142
    ._dfc_wire_104                          (_ADD124__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:270:130
    ._dfc_wire_107                          (_MUL125__dfc_wire_107)
  );
  MUL_2x1 MUL126 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:272:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_9_3152_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3170:138
    ._dfc_wire_104                          (_dup122__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:268:111
    ._dfc_wire_107                          (_MUL126__dfc_wire_107)
  );
  dup_1x2 dup127 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:273:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL125__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:271:131
    ._dfc_wire_68_105 (_dup127__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup127__dfc_wire_68_113)
  );
  ADD_2x1 ADD128 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:274:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup127__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:273:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_117_3148_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3166:146
    ._dfc_wire_100                          (_ADD128__dfc_wire_100)
  );
  MUL_2x1 MUL129 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:275:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_107_3145_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3163:146
    ._dfc_wire_104                          (_dup123__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:269:111
    ._dfc_wire_107                          (_MUL129__dfc_wire_107)
  );
  SUB_2x1 SUB130 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:276:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup127__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:273:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_27_3144_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3162:142
    ._dfc_wire_121    (_SUB130__dfc_wire_121)
  );
  dup_1x2 dup131 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:277:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST117__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:263:84
    ._dfc_wire_68_105 (_dup131__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup131__dfc_wire_68_113)
  );
  dup_1x2 dup132 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:278:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST118__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:264:84
    ._dfc_wire_68_105 (_dup132__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup132__dfc_wire_68_113)
  );
  ADD_2x1 ADD133 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:279:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup131__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:277:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_22_3143_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3161:142
    ._dfc_wire_100                          (_ADD133__dfc_wire_100)
  );
  MUL_2x1 MUL134 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:280:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_178_3142_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3160:146
    ._dfc_wire_104                          (_ADD133__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:279:130
    ._dfc_wire_107                          (_MUL134__dfc_wire_107)
  );
  MUL_2x1 MUL135 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:281:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_26_3141_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3159:142
    ._dfc_wire_104                          (_dup131__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:277:111
    ._dfc_wire_107                          (_MUL135__dfc_wire_107)
  );
  dup_1x2 dup136 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:282:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL134__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:280:131
    ._dfc_wire_68_105 (_dup136__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup136__dfc_wire_68_113)
  );
  SUB_2x1 SUB137 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:283:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup136__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:282:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_98_3140_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3158:142
    ._dfc_wire_121    (_SUB137__dfc_wire_121)
  );
  MUL_2x1 MUL138 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:284:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_62_3139_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3157:142
    ._dfc_wire_104                          (_dup132__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:278:111
    ._dfc_wire_107                          (_MUL138__dfc_wire_107)
  );
  SUB_2x1 SUB139 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:285:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup136__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:282:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_138_3138_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3156:146
    ._dfc_wire_121    (_SUB139__dfc_wire_121)
  );
  dup_1x2 dup140 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:286:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD121__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:267:130
    ._dfc_wire_68_105 (_dup140__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup140__dfc_wire_68_113)
  );
  dup_1x2 dup141 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:287:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHL11112__dfc_wire_75),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:258:89
    ._dfc_wire_68_105 (_dup141__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup141__dfc_wire_68_113)
  );
  ADD_2x1 ADD142 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:288:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup140__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:286:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_162_3137_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3155:146
    ._dfc_wire_100                          (_ADD142__dfc_wire_100)
  );
  SUB_2x1 SUB143 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:289:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup140__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:286:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_162_3136_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3154:146
    ._dfc_wire_121    (_SUB143__dfc_wire_121)
  );
  dup_1x2 dup144 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:290:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST114__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:260:84
    ._dfc_wire_68_105 (_dup144__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup144__dfc_wire_68_113)
  );
  dup_1x2 dup145 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:291:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST113__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:259:84
    ._dfc_wire_68_105 (_dup145__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup145__dfc_wire_68_113)
  );
  ADD_2x1 ADD146 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:292:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup144__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:290:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_91_3135_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3153:142
    ._dfc_wire_100                          (_ADD146__dfc_wire_100)
  );
  MUL_2x1 MUL147 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:293:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_190_3134_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3152:146
    ._dfc_wire_104                          (_ADD146__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:292:130
    ._dfc_wire_107                          (_MUL147__dfc_wire_107)
  );
  MUL_2x1 MUL148 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:294:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_9_3133_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3151:138
    ._dfc_wire_104                          (_dup145__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:291:111
    ._dfc_wire_107                          (_MUL148__dfc_wire_107)
  );
  dup_1x2 dup149 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:295:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL147__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:293:131
    ._dfc_wire_68_105 (_dup149__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup149__dfc_wire_68_113)
  );
  SUB_2x1 SUB150 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:296:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup149__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:295:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_172_3132_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3150:146
    ._dfc_wire_121    (_SUB150__dfc_wire_121)
  );
  MUL_2x1 MUL151 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:297:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_156_3131_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3149:146
    ._dfc_wire_104                          (_dup144__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:290:111
    ._dfc_wire_107                          (_MUL151__dfc_wire_107)
  );
  ADD_2x1 ADD152 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:298:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup149__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:295:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_98_3130_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3148:142
    ._dfc_wire_100                          (_ADD152__dfc_wire_100)
  );
  dup_1x2 dup153 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:299:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD128__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:274:130
    ._dfc_wire_68_105 (_dup153__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup153__dfc_wire_68_113)
  );
  dup_1x2 dup154 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:300:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB137__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:283:109
    ._dfc_wire_68_105 (_dup154__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup154__dfc_wire_68_113)
  );
  ADD_2x1 ADD155 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:301:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_51_3129_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3147:142
    .const_fix_32_0_1__0000000000000080_102 (_dup154__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:300:111
    ._dfc_wire_100                          (_ADD155__dfc_wire_100)
  );
  SUB_2x1 SUB156 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:302:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_51_3128_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3146:142
    ._dfc_wire_118    (_dup154__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:300:111
    ._dfc_wire_121    (_SUB156__dfc_wire_121)
  );
  dup_1x2 dup157 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:303:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB130__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:276:109
    ._dfc_wire_68_105 (_dup157__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup157__dfc_wire_68_113)
  );
  dup_1x2 dup158 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:304:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB139__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:285:109
    ._dfc_wire_68_105 (_dup158__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup158__dfc_wire_68_113)
  );
  ADD_2x1 ADD159 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:305:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_24_3127_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3145:142
    .const_fix_32_0_1__0000000000000080_102 (_dup158__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:304:111
    ._dfc_wire_100                          (_ADD159__dfc_wire_100)
  );
  SUB_2x1 SUB160 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:306:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_24_3126_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3144:142
    ._dfc_wire_118    (_dup158__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:304:111
    ._dfc_wire_121    (_SUB160__dfc_wire_121)
  );
  dup_1x2 dup161 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:307:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD142__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:288:130
    ._dfc_wire_68_105 (_dup161__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup161__dfc_wire_68_113)
  );
  dup_1x2 dup162 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:308:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD152__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:298:130
    ._dfc_wire_68_105 (_dup162__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup162__dfc_wire_68_113)
  );
  ADD_2x1 ADD163 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:309:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup161__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:307:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_41_3125_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3143:142
    ._dfc_wire_100                          (_ADD163__dfc_wire_100)
  );
  SUB_2x1 SUB164 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:310:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup161__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:307:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_41_3124_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3142:142
    ._dfc_wire_121    (_SUB164__dfc_wire_121)
  );
  dup_1x2 dup165 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:311:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB143__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:289:109
    ._dfc_wire_68_105 (_dup165__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup165__dfc_wire_68_113)
  );
  dup_1x2 dup166 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:312:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB150__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:296:109
    ._dfc_wire_68_105 (_dup166__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup166__dfc_wire_68_113)
  );
  ADD_2x1 ADD167 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:313:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_14_3123_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3141:142
    .const_fix_32_0_1__0000000000000080_102 (_dup166__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:312:111
    ._dfc_wire_100                          (_ADD167__dfc_wire_100)
  );
  SUB_2x1 SUB168 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:314:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_14_3122_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3140:142
    ._dfc_wire_118    (_dup166__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:312:111
    ._dfc_wire_121    (_SUB168__dfc_wire_121)
  );
  dup_1x2 dup169 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:315:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB156__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:302:109
    ._dfc_wire_68_105 (_dup169__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup169__dfc_wire_68_113)
  );
  dup_1x2 dup170 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:316:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB160__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:306:109
    ._dfc_wire_68_105 (_dup170__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup170__dfc_wire_68_113)
  );
  ADD_2x1 ADD171 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:317:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup169__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:315:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_124_3121_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3139:146
    ._dfc_wire_100                          (_ADD171__dfc_wire_100)
  );
  MUL_2x1 MUL172 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:318:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_486_3120_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3138:146
    ._dfc_wire_104                          (_ADD171__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:317:130
    ._dfc_wire_107                          (_MUL172__dfc_wire_107)
  );
  ADD_2x1 ADD173 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:319:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL172__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:318:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_636_3119_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3137:146
    ._dfc_wire_100                          (_ADD173__dfc_wire_100)
  );
  SHR8_1x1 SHR8174 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:320:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD173__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:319:130
    ._dfc_wire_216 (_SHR8174__dfc_wire_216)
  );
  SUB_2x1 SUB175 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:321:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup169__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:315:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_124_3118_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3136:146
    ._dfc_wire_121    (_SUB175__dfc_wire_121)
  );
  MUL_2x1 MUL176 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:322:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_493_3117_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3135:146
    ._dfc_wire_104                          (_SUB175__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:321:109
    ._dfc_wire_107                          (_MUL176__dfc_wire_107)
  );
  ADD_2x1 ADD177 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:323:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL176__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:322:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_624_3116_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3134:146
    ._dfc_wire_100                          (_ADD177__dfc_wire_100)
  );
  SHR8_1x1 SHR8178 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:324:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD177__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:323:130
    ._dfc_wire_216 (_SHR8178__dfc_wire_216)
  );
  dup_1x2 dup179 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:325:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD163__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:309:130
    ._dfc_wire_68_105 (_dup179__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup179__dfc_wire_68_113)
  );
  dup_1x2 dup180 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:326:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD155__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:301:130
    ._dfc_wire_68_105 (_dup180__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup180__dfc_wire_68_113)
  );
  ADD_2x1 ADD181 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:327:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_31_3115_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3133:142
    .const_fix_32_0_1__0000000000000080_102 (_dup180__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:326:111
    ._dfc_wire_100                          (_ADD181__dfc_wire_100)
  );
  SHR8_1x1 SHR8182 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:328:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD181__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:327:130
    ._dfc_wire_216 (_SHR8182__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST183 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:329:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8182__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:328:87
    ._dfc_wire_236 (_CAST183__dfc_wire_236)
  );
  dup_1x2 dup184 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:330:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD167__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:313:130
    ._dfc_wire_68_105 (_dup184__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup184__dfc_wire_68_113)
  );
  dup_1x2 dup185 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:331:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR8174__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:320:87
    ._dfc_wire_68_105 (_dup185__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup185__dfc_wire_68_113)
  );
  ADD_2x1 ADD186 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:332:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_461_3114_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3132:146
    .const_fix_32_0_1__0000000000000080_102 (_dup185__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:331:111
    ._dfc_wire_100                          (_ADD186__dfc_wire_100)
  );
  SHR8_1x1 SHR8187 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:333:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD186__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:332:130
    ._dfc_wire_216 (_SHR8187__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST188 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:334:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8187__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:333:87
    ._dfc_wire_236 (_CAST188__dfc_wire_236)
  );
  dup_1x2 dup189 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:335:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB168__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:314:109
    ._dfc_wire_68_105 (_dup189__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup189__dfc_wire_68_113)
  );
  dup_1x2 dup190 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:336:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR8178__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:324:87
    ._dfc_wire_68_105 (_dup190__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup190__dfc_wire_68_113)
  );
  ADD_2x1 ADD191 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:337:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_184_3113_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3131:146
    .const_fix_32_0_1__0000000000000080_102 (_dup190__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:336:111
    ._dfc_wire_100                          (_ADD191__dfc_wire_100)
  );
  SHR8_1x1 SHR8192 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:338:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD191__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:337:130
    ._dfc_wire_216 (_SHR8192__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST193 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:339:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8192__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:338:87
    ._dfc_wire_236 (_CAST193__dfc_wire_236)
  );
  dup_1x2 dup194 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:340:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB164__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:310:109
    ._dfc_wire_68_105 (_dup194__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup194__dfc_wire_68_113)
  );
  dup_1x2 dup195 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:341:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD159__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:305:130
    ._dfc_wire_68_105 (_dup195__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup195__dfc_wire_68_113)
  );
  ADD_2x1 ADD196 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:342:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup194__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:340:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_110_3112_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3130:146
    ._dfc_wire_100                          (_ADD196__dfc_wire_100)
  );
  SHR8_1x1 SHR8197 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:343:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD196__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:342:130
    ._dfc_wire_216 (_SHR8197__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST198 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:344:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8197__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:343:87
    ._dfc_wire_236 (_CAST198__dfc_wire_236)
  );
  SUB_2x1 SUB199 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:345:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup194__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:340:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_110_3111_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3129:146
    ._dfc_wire_121    (_SUB199__dfc_wire_121)
  );
  SHR8_1x1 SHR8200 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:346:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB199__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:345:109
    ._dfc_wire_216 (_SHR8200__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST201 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:347:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8200__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:346:87
    ._dfc_wire_236 (_CAST201__dfc_wire_236)
  );
  SUB_2x1 SUB202 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:348:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_184_3110_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3128:146
    ._dfc_wire_118    (_dup190__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:336:111
    ._dfc_wire_121    (_SUB202__dfc_wire_121)
  );
  SHR8_1x1 SHR8203 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:349:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB202__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:348:109
    ._dfc_wire_216 (_SHR8203__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST204 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:350:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8203__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:349:87
    ._dfc_wire_236 (_CAST204__dfc_wire_236)
  );
  SUB_2x1 SUB205 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:351:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_461_3109_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3127:146
    ._dfc_wire_118    (_dup185__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:331:111
    ._dfc_wire_121    (_SUB205__dfc_wire_121)
  );
  SHR8_1x1 SHR8206 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:352:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB205__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:351:109
    ._dfc_wire_216 (_SHR8206__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST207 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:353:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8206__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:352:87
    ._dfc_wire_236 (_CAST207__dfc_wire_236)
  );
  SUB_2x1 SUB208 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:354:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_31_3108_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3126:142
    ._dfc_wire_118    (_dup180__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:326:111
    ._dfc_wire_121    (_SUB208__dfc_wire_121)
  );
  SHR8_1x1 SHR8209 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:355:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB208__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:354:109
    ._dfc_wire_216 (_SHR8209__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST210 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:356:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8209__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:355:87
    ._dfc_wire_236 (_CAST210__dfc_wire_236)
  );
  CAST_1x1_16_32 CAST211 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:357:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_20__dfc_wire_45),
    ._dfc_wire_73 (_CAST211__dfc_wire_73)
  );
  SHL11_1x1 SHL11212 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:358:89
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_73 (_CAST211__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:357:84
    ._dfc_wire_75 (_SHL11212__dfc_wire_75)
  );
  CAST_1x1_16_32 CAST213 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:359:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_22__dfc_wire_45),
    ._dfc_wire_73 (_CAST213__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST214 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:360:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_18__dfc_wire_45),
    ._dfc_wire_73 (_CAST214__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST215 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:361:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_17__dfc_wire_45),
    ._dfc_wire_73 (_CAST215__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST216 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:362:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_23__dfc_wire_45),
    ._dfc_wire_73 (_CAST216__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST217 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:363:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_21__dfc_wire_45),
    ._dfc_wire_73 (_CAST217__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST218 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:364:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_19__dfc_wire_45),
    ._dfc_wire_73 (_CAST218__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST219 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:365:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_16__dfc_wire_45),
    ._dfc_wire_73 (_CAST219__dfc_wire_73)
  );
  SHL11_1x1 SHL11220 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:366:89
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_73 (_CAST219__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:365:84
    ._dfc_wire_75 (_SHL11220__dfc_wire_75)
  );
  ADD_2x1 ADD221 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:367:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_SHL11220__dfc_wire_75),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:366:89
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_97_3107_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3125:142
    ._dfc_wire_100                          (_ADD221__dfc_wire_100)
  );
  dup_1x2 dup222 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:368:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST215__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:361:84
    ._dfc_wire_68_105 (_dup222__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup222__dfc_wire_68_113)
  );
  dup_1x2 dup223 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:369:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST216__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:362:84
    ._dfc_wire_68_105 (_dup223__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup223__dfc_wire_68_113)
  );
  ADD_2x1 ADD224 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:370:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup222__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:368:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_13_3105_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3123:142
    ._dfc_wire_100                          (_ADD224__dfc_wire_100)
  );
  MUL_2x1 MUL225 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:371:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_143_3104_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3122:146
    ._dfc_wire_104                          (_ADD224__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:370:130
    ._dfc_wire_107                          (_MUL225__dfc_wire_107)
  );
  MUL_2x1 MUL226 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:372:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_66_3103_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3121:142
    ._dfc_wire_104                          (_dup222__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:368:111
    ._dfc_wire_107                          (_MUL226__dfc_wire_107)
  );
  dup_1x2 dup227 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:373:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL225__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:371:131
    ._dfc_wire_68_105 (_dup227__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup227__dfc_wire_68_113)
  );
  ADD_2x1 ADD228 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:374:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup227__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:373:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_225_3102_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3120:146
    ._dfc_wire_100                          (_ADD228__dfc_wire_100)
  );
  MUL_2x1 MUL229 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:375:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_97_3101_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3119:142
    ._dfc_wire_104                          (_dup223__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:369:111
    ._dfc_wire_107                          (_MUL229__dfc_wire_107)
  );
  SUB_2x1 SUB230 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:376:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup227__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:373:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_212_3100_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3118:146
    ._dfc_wire_121    (_SUB230__dfc_wire_121)
  );
  dup_1x2 dup231 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:377:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST217__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:363:84
    ._dfc_wire_68_105 (_dup231__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup231__dfc_wire_68_113)
  );
  dup_1x2 dup232 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:378:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST218__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:364:84
    ._dfc_wire_68_105 (_dup232__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup232__dfc_wire_68_113)
  );
  ADD_2x1 ADD233 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:379:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_52_3099_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3117:142
    .const_fix_32_0_1__0000000000000080_102 (_dup232__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:378:111
    ._dfc_wire_100                          (_ADD233__dfc_wire_100)
  );
  MUL_2x1 MUL234 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:380:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_256_3098_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3116:146
    ._dfc_wire_104                          (_ADD233__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:379:130
    ._dfc_wire_107                          (_MUL234__dfc_wire_107)
  );
  MUL_2x1 MUL235 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:381:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_50_3097_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3115:142
    ._dfc_wire_104                          (_dup231__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:377:111
    ._dfc_wire_107                          (_MUL235__dfc_wire_107)
  );
  dup_1x2 dup236 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:382:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL234__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:380:131
    ._dfc_wire_68_105 (_dup236__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup236__dfc_wire_68_113)
  );
  SUB_2x1 SUB237 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:383:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup236__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:382:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_146_3096_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3114:146
    ._dfc_wire_121    (_SUB237__dfc_wire_121)
  );
  MUL_2x1 MUL238 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:384:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_160_3095_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3113:146
    ._dfc_wire_104                          (_dup232__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:378:111
    ._dfc_wire_107                          (_MUL238__dfc_wire_107)
  );
  SUB_2x1 SUB239 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:385:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup236__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:382:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_143_3093_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3111:146
    ._dfc_wire_121    (_SUB239__dfc_wire_121)
  );
  dup_1x2 dup240 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:386:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD221__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:367:130
    ._dfc_wire_68_105 (_dup240__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup240__dfc_wire_68_113)
  );
  dup_1x2 dup241 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:387:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHL11212__dfc_wire_75),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:358:89
    ._dfc_wire_68_105 (_dup241__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup241__dfc_wire_68_113)
  );
  ADD_2x1 ADD242 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:388:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_53_3092_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3110:142
    .const_fix_32_0_1__0000000000000080_102 (_dup241__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:387:111
    ._dfc_wire_100                          (_ADD242__dfc_wire_100)
  );
  SUB_2x1 SUB243 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:389:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_53_3091_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3109:142
    ._dfc_wire_118    (_dup241__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:387:111
    ._dfc_wire_121    (_SUB243__dfc_wire_121)
  );
  dup_1x2 dup244 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:390:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST214__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:360:84
    ._dfc_wire_68_105 (_dup244__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup244__dfc_wire_68_113)
  );
  dup_1x2 dup245 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:391:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST213__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:359:84
    ._dfc_wire_68_105 (_dup245__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup245__dfc_wire_68_113)
  );
  ADD_2x1 ADD246 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:392:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup244__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:390:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_15_3089_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3107:142
    ._dfc_wire_100                          (_ADD246__dfc_wire_100)
  );
  MUL_2x1 MUL247 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:393:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_83_3088_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3106:142
    ._dfc_wire_104                          (_ADD246__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:392:130
    ._dfc_wire_107                          (_MUL247__dfc_wire_107)
  );
  MUL_2x1 MUL248 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:394:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_39_3087_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3105:142
    ._dfc_wire_104                          (_dup245__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:391:111
    ._dfc_wire_107                          (_MUL248__dfc_wire_107)
  );
  dup_1x2 dup249 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:395:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL247__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:393:131
    ._dfc_wire_68_105 (_dup249__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup249__dfc_wire_68_113)
  );
  SUB_2x1 SUB250 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:396:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup249__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:395:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_110_3085_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3103:146
    ._dfc_wire_121    (_SUB250__dfc_wire_121)
  );
  MUL_2x1 MUL251 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:397:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_110_3084_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3102:146
    ._dfc_wire_104                          (_dup244__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:390:111
    ._dfc_wire_107                          (_MUL251__dfc_wire_107)
  );
  ADD_2x1 ADD252 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:398:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup249__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:395:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_33_3082_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3100:142
    ._dfc_wire_100                          (_ADD252__dfc_wire_100)
  );
  dup_1x2 dup253 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:399:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD228__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:374:130
    ._dfc_wire_68_105 (_dup253__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup253__dfc_wire_68_113)
  );
  dup_1x2 dup254 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:400:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB237__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:383:109
    ._dfc_wire_68_105 (_dup254__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup254__dfc_wire_68_113)
  );
  ADD_2x1 ADD255 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:401:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_37_3080_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3098:142
    .const_fix_32_0_1__0000000000000080_102 (_dup254__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:400:111
    ._dfc_wire_100                          (_ADD255__dfc_wire_100)
  );
  SUB_2x1 SUB256 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:402:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_37_3079_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3097:142
    ._dfc_wire_118    (_dup254__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:400:111
    ._dfc_wire_121    (_SUB256__dfc_wire_121)
  );
  dup_1x2 dup257 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:403:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB230__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:376:109
    ._dfc_wire_68_105 (_dup257__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup257__dfc_wire_68_113)
  );
  dup_1x2 dup258 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:404:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB239__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:385:109
    ._dfc_wire_68_105 (_dup258__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup258__dfc_wire_68_113)
  );
  ADD_2x1 ADD259 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:405:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_28_3077_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3095:142
    .const_fix_32_0_1__0000000000000080_102 (_dup258__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:404:111
    ._dfc_wire_100                          (_ADD259__dfc_wire_100)
  );
  SUB_2x1 SUB260 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:406:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_28_3076_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3094:142
    ._dfc_wire_118    (_dup258__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:404:111
    ._dfc_wire_121    (_SUB260__dfc_wire_121)
  );
  dup_1x2 dup261 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:407:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD242__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:388:130
    ._dfc_wire_68_105 (_dup261__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup261__dfc_wire_68_113)
  );
  dup_1x2 dup262 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:408:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD252__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:398:130
    ._dfc_wire_68_105 (_dup262__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup262__dfc_wire_68_113)
  );
  ADD_2x1 ADD263 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:409:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup261__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:407:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_47_3072_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3090:142
    ._dfc_wire_100                          (_ADD263__dfc_wire_100)
  );
  SUB_2x1 SUB264 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:410:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup261__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:407:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_47_3070_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3088:142
    ._dfc_wire_121    (_SUB264__dfc_wire_121)
  );
  dup_1x2 dup265 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:411:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB243__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:389:109
    ._dfc_wire_68_105 (_dup265__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup265__dfc_wire_68_113)
  );
  dup_1x2 dup266 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:412:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB250__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:396:109
    ._dfc_wire_68_105 (_dup266__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup266__dfc_wire_68_113)
  );
  ADD_2x1 ADD267 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:413:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup265__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:411:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_51_3064_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3082:142
    ._dfc_wire_100                          (_ADD267__dfc_wire_100)
  );
  SUB_2x1 SUB268 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:414:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup265__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:411:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_51_3061_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3079:142
    ._dfc_wire_121    (_SUB268__dfc_wire_121)
  );
  dup_1x2 dup269 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:415:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB256__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:402:109
    ._dfc_wire_68_105 (_dup269__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup269__dfc_wire_68_113)
  );
  dup_1x2 dup270 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:416:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB260__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:406:109
    ._dfc_wire_68_105 (_dup270__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup270__dfc_wire_68_113)
  );
  ADD_2x1 ADD271 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:417:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup269__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:415:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_31_3051_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3069:142
    ._dfc_wire_100                          (_ADD271__dfc_wire_100)
  );
  MUL_2x1 MUL272 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:418:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_574_3049_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3067:146
    ._dfc_wire_104                          (_ADD271__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:417:130
    ._dfc_wire_107                          (_MUL272__dfc_wire_107)
  );
  ADD_2x1 ADD273 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:419:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL272__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:418:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_717_3047_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3065:146
    ._dfc_wire_100                          (_ADD273__dfc_wire_100)
  );
  SHR8_1x1 SHR8274 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:420:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD273__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:419:130
    ._dfc_wire_216 (_SHR8274__dfc_wire_216)
  );
  SUB_2x1 SUB275 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:421:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup269__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:415:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_31_3045_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3063:142
    ._dfc_wire_121    (_SUB275__dfc_wire_121)
  );
  MUL_2x1 MUL276 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:422:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_634_3041_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3059:146
    ._dfc_wire_104                          (_SUB275__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:421:109
    ._dfc_wire_107                          (_MUL276__dfc_wire_107)
  );
  ADD_2x1 ADD277 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:423:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL276__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:422:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_778_3037_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3055:146
    ._dfc_wire_100                          (_ADD277__dfc_wire_100)
  );
  SHR8_1x1 SHR8278 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:424:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD277__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:423:130
    ._dfc_wire_216 (_SHR8278__dfc_wire_216)
  );
  dup_1x2 dup279 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:425:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD263__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:409:130
    ._dfc_wire_68_105 (_dup279__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup279__dfc_wire_68_113)
  );
  dup_1x2 dup280 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:426:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD255__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:401:130
    ._dfc_wire_68_105 (_dup280__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup280__dfc_wire_68_113)
  );
  ADD_2x1 ADD281 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:427:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_94_3029_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3047:142
    .const_fix_32_0_1__0000000000000080_102 (_dup280__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:426:111
    ._dfc_wire_100                          (_ADD281__dfc_wire_100)
  );
  SHR8_1x1 SHR8282 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:428:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD281__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:427:130
    ._dfc_wire_216 (_SHR8282__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST283 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:429:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8282__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:428:87
    ._dfc_wire_236 (_CAST283__dfc_wire_236)
  );
  dup_1x2 dup284 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:430:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD267__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:413:130
    ._dfc_wire_68_105 (_dup284__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup284__dfc_wire_68_113)
  );
  dup_1x2 dup285 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:431:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR8274__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:420:87
    ._dfc_wire_68_105 (_dup285__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup285__dfc_wire_68_113)
  );
  ADD_2x1 ADD286 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:432:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_399_3019_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3037:146
    .const_fix_32_0_1__0000000000000080_102 (_dup285__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:431:111
    ._dfc_wire_100                          (_ADD286__dfc_wire_100)
  );
  SHR8_1x1 SHR8287 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:433:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD286__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:432:130
    ._dfc_wire_216 (_SHR8287__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST288 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:434:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8287__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:433:87
    ._dfc_wire_236 (_CAST288__dfc_wire_236)
  );
  dup_1x2 dup289 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:435:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB268__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:414:109
    ._dfc_wire_68_105 (_dup289__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup289__dfc_wire_68_113)
  );
  dup_1x2 dup290 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:436:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR8278__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:424:87
    ._dfc_wire_68_105 (_dup290__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup290__dfc_wire_68_113)
  );
  ADD_2x1 ADD291 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:437:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_480_3011_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3029:146
    .const_fix_32_0_1__0000000000000080_102 (_dup290__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:436:111
    ._dfc_wire_100                          (_ADD291__dfc_wire_100)
  );
  SHR8_1x1 SHR8292 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:438:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD291__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:437:130
    ._dfc_wire_216 (_SHR8292__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST293 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:439:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8292__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:438:87
    ._dfc_wire_236 (_CAST293__dfc_wire_236)
  );
  dup_1x2 dup294 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:440:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB264__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:410:109
    ._dfc_wire_68_105 (_dup294__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup294__dfc_wire_68_113)
  );
  dup_1x2 dup295 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:441:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD259__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:405:130
    ._dfc_wire_68_105 (_dup295__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup295__dfc_wire_68_113)
  );
  ADD_2x1 ADD296 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:442:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_90_2997_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3015:142
    .const_fix_32_0_1__0000000000000080_102 (_dup295__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:441:111
    ._dfc_wire_100                          (_ADD296__dfc_wire_100)
  );
  SHR8_1x1 SHR8297 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:443:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD296__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:442:130
    ._dfc_wire_216 (_SHR8297__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST298 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:444:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8297__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:443:87
    ._dfc_wire_236 (_CAST298__dfc_wire_236)
  );
  SUB_2x1 SUB299 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:445:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_90_3212_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3230:142
    ._dfc_wire_118    (_dup295__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:441:111
    ._dfc_wire_121    (_SUB299__dfc_wire_121)
  );
  SHR8_1x1 SHR8300 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:446:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB299__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:445:109
    ._dfc_wire_216 (_SHR8300__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST301 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:447:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8300__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:446:87
    ._dfc_wire_236 (_CAST301__dfc_wire_236)
  );
  SUB_2x1 SUB302 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:448:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_480_2993_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3011:146
    ._dfc_wire_118    (_dup290__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:436:111
    ._dfc_wire_121    (_SUB302__dfc_wire_121)
  );
  SHR8_1x1 SHR8303 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:449:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB302__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:448:109
    ._dfc_wire_216 (_SHR8303__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST304 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:450:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8303__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:449:87
    ._dfc_wire_236 (_CAST304__dfc_wire_236)
  );
  SUB_2x1 SUB305 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:451:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_399_2988_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3006:146
    ._dfc_wire_118    (_dup285__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:431:111
    ._dfc_wire_121    (_SUB305__dfc_wire_121)
  );
  SHR8_1x1 SHR8306 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:452:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB305__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:451:109
    ._dfc_wire_216 (_SHR8306__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST307 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:453:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8306__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:452:87
    ._dfc_wire_236 (_CAST307__dfc_wire_236)
  );
  SUB_2x1 SUB308 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:454:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_94_2984_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3002:142
    ._dfc_wire_118    (_dup280__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:426:111
    ._dfc_wire_121    (_SUB308__dfc_wire_121)
  );
  SHR8_1x1 SHR8309 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:455:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB308__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:454:109
    ._dfc_wire_216 (_SHR8309__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST310 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:456:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8309__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:455:87
    ._dfc_wire_236 (_CAST310__dfc_wire_236)
  );
  CAST_1x1_16_32 CAST311 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:457:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_28__dfc_wire_45),
    ._dfc_wire_73 (_CAST311__dfc_wire_73)
  );
  SHL11_1x1 SHL11312 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:458:89
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_73 (_CAST311__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:457:84
    ._dfc_wire_75 (_SHL11312__dfc_wire_75)
  );
  CAST_1x1_16_32 CAST313 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:459:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_30__dfc_wire_45),
    ._dfc_wire_73 (_CAST313__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST314 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:460:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_26__dfc_wire_45),
    ._dfc_wire_73 (_CAST314__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST315 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:461:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_25__dfc_wire_45),
    ._dfc_wire_73 (_CAST315__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST316 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:462:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_31__dfc_wire_45),
    ._dfc_wire_73 (_CAST316__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST317 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:463:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_29__dfc_wire_45),
    ._dfc_wire_73 (_CAST317__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST318 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:464:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_27__dfc_wire_45),
    ._dfc_wire_73 (_CAST318__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST319 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:465:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_24__dfc_wire_45),
    ._dfc_wire_73 (_CAST319__dfc_wire_73)
  );
  SHL11_1x1 SHL11320 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:466:89
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_73 (_CAST319__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:465:84
    ._dfc_wire_75 (_SHL11320__dfc_wire_75)
  );
  ADD_2x1 ADD321 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:467:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_SHL11320__dfc_wire_75),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:466:89
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_122_2977_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2995:146
    ._dfc_wire_100                          (_ADD321__dfc_wire_100)
  );
  dup_1x2 dup322 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:468:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST315__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:461:84
    ._dfc_wire_68_105 (_dup322__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup322__dfc_wire_68_113)
  );
  dup_1x2 dup323 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:469:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST316__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:462:84
    ._dfc_wire_68_105 (_dup323__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup323__dfc_wire_68_113)
  );
  ADD_2x1 ADD324 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:470:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_54_2976_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2994:142
    .const_fix_32_0_1__0000000000000080_102 (_dup323__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:469:111
    ._dfc_wire_100                          (_ADD324__dfc_wire_100)
  );
  MUL_2x1 MUL325 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:471:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_113_2975_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2993:146
    ._dfc_wire_104                          (_ADD324__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:470:130
    ._dfc_wire_107                          (_MUL325__dfc_wire_107)
  );
  MUL_2x1 MUL326 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:472:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_44_2974_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2992:142
    ._dfc_wire_104                          (_dup322__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:468:111
    ._dfc_wire_107                          (_MUL326__dfc_wire_107)
  );
  dup_1x2 dup327 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:473:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL325__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:471:131
    ._dfc_wire_68_105 (_dup327__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup327__dfc_wire_68_113)
  );
  ADD_2x1 ADD328 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:474:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup327__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:473:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_60_2973_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2991:142
    ._dfc_wire_100                          (_ADD328__dfc_wire_100)
  );
  MUL_2x1 MUL329 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:475:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_142_2972_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2990:146
    ._dfc_wire_104                          (_dup323__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:469:111
    ._dfc_wire_107                          (_MUL329__dfc_wire_107)
  );
  SUB_2x1 SUB330 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:476:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup327__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:473:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_39_2971_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2989:142
    ._dfc_wire_121    (_SUB330__dfc_wire_121)
  );
  dup_1x2 dup331 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:477:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST317__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:463:84
    ._dfc_wire_68_105 (_dup331__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup331__dfc_wire_68_113)
  );
  dup_1x2 dup332 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:478:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST318__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:464:84
    ._dfc_wire_68_105 (_dup332__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup332__dfc_wire_68_113)
  );
  ADD_2x1 ADD333 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:479:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup331__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:477:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_76_2970_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2988:142
    ._dfc_wire_100                          (_ADD333__dfc_wire_100)
  );
  MUL_2x1 MUL334 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:480:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_199_2969_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2987:146
    ._dfc_wire_104                          (_ADD333__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:479:130
    ._dfc_wire_107                          (_MUL334__dfc_wire_107)
  );
  MUL_2x1 MUL335 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:481:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_43_2968_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2986:142
    ._dfc_wire_104                          (_dup331__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:477:111
    ._dfc_wire_107                          (_MUL335__dfc_wire_107)
  );
  dup_1x2 dup336 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:482:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL334__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:480:131
    ._dfc_wire_68_105 (_dup336__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup336__dfc_wire_68_113)
  );
  SUB_2x1 SUB337 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:483:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup336__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:482:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_94_2967_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2985:142
    ._dfc_wire_121    (_SUB337__dfc_wire_121)
  );
  MUL_2x1 MUL338 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:484:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_25_2966_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2984:142
    ._dfc_wire_104                          (_dup332__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:478:111
    ._dfc_wire_107                          (_MUL338__dfc_wire_107)
  );
  SUB_2x1 SUB339 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:485:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup336__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:482:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_186_2965_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2983:146
    ._dfc_wire_121    (_SUB339__dfc_wire_121)
  );
  dup_1x2 dup340 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:486:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD321__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:467:130
    ._dfc_wire_68_105 (_dup340__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup340__dfc_wire_68_113)
  );
  dup_1x2 dup341 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:487:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHL11312__dfc_wire_75),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:458:89
    ._dfc_wire_68_105 (_dup341__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup341__dfc_wire_68_113)
  );
  ADD_2x1 ADD342 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:488:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_12_2964_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2982:142
    .const_fix_32_0_1__0000000000000080_102 (_dup341__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:487:111
    ._dfc_wire_100                          (_ADD342__dfc_wire_100)
  );
  SUB_2x1 SUB343 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:489:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_12_2963_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2981:142
    ._dfc_wire_118    (_dup341__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:487:111
    ._dfc_wire_121    (_SUB343__dfc_wire_121)
  );
  dup_1x2 dup344 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:490:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST314__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:460:84
    ._dfc_wire_68_105 (_dup344__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup344__dfc_wire_68_113)
  );
  dup_1x2 dup345 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:491:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST313__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:459:84
    ._dfc_wire_68_105 (_dup345__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup345__dfc_wire_68_113)
  );
  ADD_2x1 ADD346 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:492:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_72_2962_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2980:142
    .const_fix_32_0_1__0000000000000080_102 (_dup345__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:491:111
    ._dfc_wire_100                          (_ADD346__dfc_wire_100)
  );
  MUL_2x1 MUL347 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:493:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_136_2961_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2979:146
    ._dfc_wire_104                          (_ADD346__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:492:130
    ._dfc_wire_107                          (_MUL347__dfc_wire_107)
  );
  MUL_2x1 MUL348 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:494:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_44_2960_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2978:142
    ._dfc_wire_104                          (_dup345__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:491:111
    ._dfc_wire_107                          (_MUL348__dfc_wire_107)
  );
  dup_1x2 dup349 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:495:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL347__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:493:131
    ._dfc_wire_68_105 (_dup349__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup349__dfc_wire_68_113)
  );
  SUB_2x1 SUB350 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:496:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup349__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:495:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_155_2959_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2977:146
    ._dfc_wire_121    (_SUB350__dfc_wire_121)
  );
  MUL_2x1 MUL351 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:497:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_28_2958_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2976:142
    ._dfc_wire_104                          (_dup344__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:490:111
    ._dfc_wire_107                          (_MUL351__dfc_wire_107)
  );
  ADD_2x1 ADD352 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:498:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup349__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:495:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_253_2957_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2975:146
    ._dfc_wire_100                          (_ADD352__dfc_wire_100)
  );
  dup_1x2 dup353 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:499:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD328__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:474:130
    ._dfc_wire_68_105 (_dup353__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup353__dfc_wire_68_113)
  );
  dup_1x2 dup354 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:500:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB337__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:483:109
    ._dfc_wire_68_105 (_dup354__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup354__dfc_wire_68_113)
  );
  ADD_2x1 ADD355 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:501:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_15_2956_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2974:142
    .const_fix_32_0_1__0000000000000080_102 (_dup354__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:500:111
    ._dfc_wire_100                          (_ADD355__dfc_wire_100)
  );
  SUB_2x1 SUB356 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:502:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_15_2955_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2973:142
    ._dfc_wire_118    (_dup354__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:500:111
    ._dfc_wire_121    (_SUB356__dfc_wire_121)
  );
  dup_1x2 dup357 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:503:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB330__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:476:109
    ._dfc_wire_68_105 (_dup357__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup357__dfc_wire_68_113)
  );
  dup_1x2 dup358 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:504:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB339__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:485:109
    ._dfc_wire_68_105 (_dup358__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup358__dfc_wire_68_113)
  );
  ADD_2x1 ADD359 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:505:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_16_2954_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2972:142
    .const_fix_32_0_1__0000000000000080_102 (_dup358__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:504:111
    ._dfc_wire_100                          (_ADD359__dfc_wire_100)
  );
  SUB_2x1 SUB360 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:506:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_16_2953_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2971:142
    ._dfc_wire_118    (_dup358__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:504:111
    ._dfc_wire_121    (_SUB360__dfc_wire_121)
  );
  dup_1x2 dup361 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:507:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD342__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:488:130
    ._dfc_wire_68_105 (_dup361__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup361__dfc_wire_68_113)
  );
  dup_1x2 dup362 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:508:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD352__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:498:130
    ._dfc_wire_68_105 (_dup362__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup362__dfc_wire_68_113)
  );
  ADD_2x1 ADD363 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:509:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_14_2952_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2970:142
    .const_fix_32_0_1__0000000000000080_102 (_dup362__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:508:111
    ._dfc_wire_100                          (_ADD363__dfc_wire_100)
  );
  SUB_2x1 SUB364 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:510:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_14_2951_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2969:142
    ._dfc_wire_118    (_dup362__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:508:111
    ._dfc_wire_121    (_SUB364__dfc_wire_121)
  );
  dup_1x2 dup365 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:511:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB343__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:489:109
    ._dfc_wire_68_105 (_dup365__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup365__dfc_wire_68_113)
  );
  dup_1x2 dup366 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:512:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB350__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:496:109
    ._dfc_wire_68_105 (_dup366__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup366__dfc_wire_68_113)
  );
  ADD_2x1 ADD367 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:513:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_87_2950_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2968:142
    .const_fix_32_0_1__0000000000000080_102 (_dup366__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:512:111
    ._dfc_wire_100                          (_ADD367__dfc_wire_100)
  );
  SUB_2x1 SUB368 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:514:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_87_2949_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2967:142
    ._dfc_wire_118    (_dup366__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:512:111
    ._dfc_wire_121    (_SUB368__dfc_wire_121)
  );
  dup_1x2 dup369 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:515:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB356__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:502:109
    ._dfc_wire_68_105 (_dup369__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup369__dfc_wire_68_113)
  );
  dup_1x2 dup370 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:516:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB360__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:506:109
    ._dfc_wire_68_105 (_dup370__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup370__dfc_wire_68_113)
  );
  ADD_2x1 ADD371 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:517:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup369__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:515:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_46_2948_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2966:142
    ._dfc_wire_100                          (_ADD371__dfc_wire_100)
  );
  MUL_2x1 MUL372 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:518:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_482_2947_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2965:146
    ._dfc_wire_104                          (_ADD371__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:517:130
    ._dfc_wire_107                          (_MUL372__dfc_wire_107)
  );
  ADD_2x1 ADD373 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:519:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL372__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:518:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_625_2946_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2964:146
    ._dfc_wire_100                          (_ADD373__dfc_wire_100)
  );
  SHR8_1x1 SHR8374 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:520:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD373__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:519:130
    ._dfc_wire_216 (_SHR8374__dfc_wire_216)
  );
  SUB_2x1 SUB375 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:521:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup369__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:515:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_46_2945_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2963:142
    ._dfc_wire_121    (_SUB375__dfc_wire_121)
  );
  MUL_2x1 MUL376 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:522:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_456_2944_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2962:146
    ._dfc_wire_104                          (_SUB375__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:521:109
    ._dfc_wire_107                          (_MUL376__dfc_wire_107)
  );
  ADD_2x1 ADD377 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:523:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL376__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:522:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_609_2943_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2961:146
    ._dfc_wire_100                          (_ADD377__dfc_wire_100)
  );
  SHR8_1x1 SHR8378 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:524:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD377__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:523:130
    ._dfc_wire_216 (_SHR8378__dfc_wire_216)
  );
  dup_1x2 dup379 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:525:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD363__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:509:130
    ._dfc_wire_68_105 (_dup379__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup379__dfc_wire_68_113)
  );
  dup_1x2 dup380 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:526:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD355__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:501:130
    ._dfc_wire_68_105 (_dup380__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup380__dfc_wire_68_113)
  );
  ADD_2x1 ADD381 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:527:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup379__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:525:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_55_2942_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2960:142
    ._dfc_wire_100                          (_ADD381__dfc_wire_100)
  );
  SHR8_1x1 SHR8382 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:528:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD381__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:527:130
    ._dfc_wire_216 (_SHR8382__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST383 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:529:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8382__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:528:87
    ._dfc_wire_236 (_CAST383__dfc_wire_236)
  );
  dup_1x2 dup384 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:530:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD367__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:513:130
    ._dfc_wire_68_105 (_dup384__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup384__dfc_wire_68_113)
  );
  dup_1x2 dup385 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:531:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR8374__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:520:87
    ._dfc_wire_68_105 (_dup385__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup385__dfc_wire_68_113)
  );
  ADD_2x1 ADD386 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:532:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_270_3094_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3112:146
    .const_fix_32_0_1__0000000000000080_102 (_dup385__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:531:111
    ._dfc_wire_100                          (_ADD386__dfc_wire_100)
  );
  SHR8_1x1 SHR8387 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:533:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD386__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:532:130
    ._dfc_wire_216 (_SHR8387__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST388 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:534:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8387__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:533:87
    ._dfc_wire_236 (_CAST388__dfc_wire_236)
  );
  dup_1x2 dup389 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:535:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB368__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:514:109
    ._dfc_wire_68_105 (_dup389__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup389__dfc_wire_68_113)
  );
  dup_1x2 dup390 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:536:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR8378__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:524:87
    ._dfc_wire_68_105 (_dup390__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup390__dfc_wire_68_113)
  );
  ADD_2x1 ADD391 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:537:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_216_3090_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3108:146
    .const_fix_32_0_1__0000000000000080_102 (_dup390__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:536:111
    ._dfc_wire_100                          (_ADD391__dfc_wire_100)
  );
  SHR8_1x1 SHR8392 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:538:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD391__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:537:130
    ._dfc_wire_216 (_SHR8392__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST393 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:539:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8392__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:538:87
    ._dfc_wire_236 (_CAST393__dfc_wire_236)
  );
  dup_1x2 dup394 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:540:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB364__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:510:109
    ._dfc_wire_68_105 (_dup394__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup394__dfc_wire_68_113)
  );
  dup_1x2 dup395 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:541:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD359__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:505:130
    ._dfc_wire_68_105 (_dup395__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup395__dfc_wire_68_113)
  );
  ADD_2x1 ADD396 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:542:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_17_3086_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3104:142
    .const_fix_32_0_1__0000000000000080_102 (_dup395__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:541:111
    ._dfc_wire_100                          (_ADD396__dfc_wire_100)
  );
  SHR8_1x1 SHR8397 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:543:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD396__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:542:130
    ._dfc_wire_216 (_SHR8397__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST398 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:544:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8397__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:543:87
    ._dfc_wire_236 (_CAST398__dfc_wire_236)
  );
  SUB_2x1 SUB399 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:545:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_17_3083_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3101:142
    ._dfc_wire_118    (_dup395__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:541:111
    ._dfc_wire_121    (_SUB399__dfc_wire_121)
  );
  SHR8_1x1 SHR8400 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:546:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB399__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:545:109
    ._dfc_wire_216 (_SHR8400__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST401 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:547:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8400__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:546:87
    ._dfc_wire_236 (_CAST401__dfc_wire_236)
  );
  SUB_2x1 SUB402 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:548:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_216_3081_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3099:146
    ._dfc_wire_118    (_dup390__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:536:111
    ._dfc_wire_121    (_SUB402__dfc_wire_121)
  );
  SHR8_1x1 SHR8403 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:549:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB402__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:548:109
    ._dfc_wire_216 (_SHR8403__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST404 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:550:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8403__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:549:87
    ._dfc_wire_236 (_CAST404__dfc_wire_236)
  );
  SUB_2x1 SUB405 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:551:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_270_2941_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2959:146
    ._dfc_wire_118    (_dup385__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:531:111
    ._dfc_wire_121    (_SUB405__dfc_wire_121)
  );
  SHR8_1x1 SHR8406 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:552:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB405__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:551:109
    ._dfc_wire_216 (_SHR8406__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST407 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:553:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8406__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:552:87
    ._dfc_wire_236 (_CAST407__dfc_wire_236)
  );
  SUB_2x1 SUB408 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:554:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup379__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:525:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_55_2940_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2958:142
    ._dfc_wire_121    (_SUB408__dfc_wire_121)
  );
  SHR8_1x1 SHR8409 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:555:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB408__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:554:109
    ._dfc_wire_216 (_SHR8409__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST410 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:556:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8409__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:555:87
    ._dfc_wire_236 (_CAST410__dfc_wire_236)
  );
  CAST_1x1_16_32 CAST411 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:557:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_36__dfc_wire_45),
    ._dfc_wire_73 (_CAST411__dfc_wire_73)
  );
  SHL11_1x1 SHL11412 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:558:89
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_73 (_CAST411__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:557:84
    ._dfc_wire_75 (_SHL11412__dfc_wire_75)
  );
  CAST_1x1_16_32 CAST413 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:559:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_38__dfc_wire_45),
    ._dfc_wire_73 (_CAST413__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST414 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:560:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_34__dfc_wire_45),
    ._dfc_wire_73 (_CAST414__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST415 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:561:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_33__dfc_wire_45),
    ._dfc_wire_73 (_CAST415__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST416 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:562:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_39__dfc_wire_45),
    ._dfc_wire_73 (_CAST416__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST417 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:563:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_37__dfc_wire_45),
    ._dfc_wire_73 (_CAST417__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST418 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:564:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_35__dfc_wire_45),
    ._dfc_wire_73 (_CAST418__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST419 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:565:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_32__dfc_wire_45),
    ._dfc_wire_73 (_CAST419__dfc_wire_73)
  );
  SHL11_1x1 SHL11420 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:566:89
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_73 (_CAST419__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:565:84
    ._dfc_wire_75 (_SHL11420__dfc_wire_75)
  );
  ADD_2x1 ADD421 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:567:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_SHL11420__dfc_wire_75),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:566:89
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_166_2934_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2952:146
    ._dfc_wire_100                          (_ADD421__dfc_wire_100)
  );
  dup_1x2 dup422 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:568:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST415__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:561:84
    ._dfc_wire_68_105 (_dup422__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup422__dfc_wire_68_113)
  );
  dup_1x2 dup423 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:569:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST416__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:562:84
    ._dfc_wire_68_105 (_dup423__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup423__dfc_wire_68_113)
  );
  ADD_2x1 ADD424 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:570:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup422__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:568:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_30_2932_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2950:142
    ._dfc_wire_100                          (_ADD424__dfc_wire_100)
  );
  MUL_2x1 MUL425 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:571:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_91_2931_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2949:142
    ._dfc_wire_104                          (_ADD424__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:570:130
    ._dfc_wire_107                          (_MUL425__dfc_wire_107)
  );
  MUL_2x1 MUL426 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:572:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_7_2930_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2948:138
    ._dfc_wire_104                          (_dup422__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:568:111
    ._dfc_wire_107                          (_MUL426__dfc_wire_107)
  );
  dup_1x2 dup427 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:573:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL425__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:571:131
    ._dfc_wire_68_105 (_dup427__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup427__dfc_wire_68_113)
  );
  ADD_2x1 ADD428 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:574:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup427__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:573:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_31_2929_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2947:142
    ._dfc_wire_100                          (_ADD428__dfc_wire_100)
  );
  MUL_2x1 MUL429 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:575:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_21_2928_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2946:142
    ._dfc_wire_104                          (_dup423__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:569:111
    ._dfc_wire_107                          (_MUL429__dfc_wire_107)
  );
  SUB_2x1 SUB430 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:576:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup427__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:573:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_89_2927_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2945:142
    ._dfc_wire_121    (_SUB430__dfc_wire_121)
  );
  dup_1x2 dup431 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:577:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST417__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:563:84
    ._dfc_wire_68_105 (_dup431__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup431__dfc_wire_68_113)
  );
  dup_1x2 dup432 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:578:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST418__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:564:84
    ._dfc_wire_68_105 (_dup432__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup432__dfc_wire_68_113)
  );
  ADD_2x1 ADD433 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:579:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_11_2926_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2944:142
    .const_fix_32_0_1__0000000000000080_102 (_dup432__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:578:111
    ._dfc_wire_100                          (_ADD433__dfc_wire_100)
  );
  MUL_2x1 MUL434 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:580:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_114_2925_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2943:146
    ._dfc_wire_104                          (_ADD433__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:579:130
    ._dfc_wire_107                          (_MUL434__dfc_wire_107)
  );
  MUL_2x1 MUL435 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:581:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_10_2924_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2942:142
    ._dfc_wire_104                          (_dup431__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:577:111
    ._dfc_wire_107                          (_MUL435__dfc_wire_107)
  );
  dup_1x2 dup436 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:582:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL434__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:580:131
    ._dfc_wire_68_105 (_dup436__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup436__dfc_wire_68_113)
  );
  SUB_2x1 SUB437 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:583:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup436__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:582:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_150_2923_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2941:146
    ._dfc_wire_121    (_SUB437__dfc_wire_121)
  );
  MUL_2x1 MUL438 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:584:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_79_2922_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2940:142
    ._dfc_wire_104                          (_dup432__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:578:111
    ._dfc_wire_107                          (_MUL438__dfc_wire_107)
  );
  SUB_2x1 SUB439 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:585:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup436__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:582:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_166_2921_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2939:146
    ._dfc_wire_121    (_SUB439__dfc_wire_121)
  );
  dup_1x2 dup440 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:586:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD421__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:567:130
    ._dfc_wire_68_105 (_dup440__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup440__dfc_wire_68_113)
  );
  dup_1x2 dup441 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:587:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHL11412__dfc_wire_75),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:558:89
    ._dfc_wire_68_105 (_dup441__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup441__dfc_wire_68_113)
  );
  ADD_2x1 ADD442 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:588:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup440__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:586:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_4_2920_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2938:138
    ._dfc_wire_100                          (_ADD442__dfc_wire_100)
  );
  SUB_2x1 SUB443 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:589:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup440__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:586:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_4_2919_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2937:138
    ._dfc_wire_121    (_SUB443__dfc_wire_121)
  );
  dup_1x2 dup444 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:590:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST414__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:560:84
    ._dfc_wire_68_105 (_dup444__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup444__dfc_wire_68_113)
  );
  dup_1x2 dup445 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:591:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST413__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:559:84
    ._dfc_wire_68_105 (_dup445__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup445__dfc_wire_68_113)
  );
  ADD_2x1 ADD446 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:592:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_66_2918_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2936:142
    .const_fix_32_0_1__0000000000000080_102 (_dup445__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:591:111
    ._dfc_wire_100                          (_ADD446__dfc_wire_100)
  );
  MUL_2x1 MUL447 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:593:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_131_2917_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2935:146
    ._dfc_wire_104                          (_ADD446__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:592:130
    ._dfc_wire_107                          (_MUL447__dfc_wire_107)
  );
  MUL_2x1 MUL448 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:594:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_81_2916_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2934:142
    ._dfc_wire_104                          (_dup445__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:591:111
    ._dfc_wire_107                          (_MUL448__dfc_wire_107)
  );
  dup_1x2 dup449 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:595:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL447__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:593:131
    ._dfc_wire_68_105 (_dup449__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup449__dfc_wire_68_113)
  );
  SUB_2x1 SUB450 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:596:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup449__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:595:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_76_2915_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2933:142
    ._dfc_wire_121    (_SUB450__dfc_wire_121)
  );
  MUL_2x1 MUL451 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:597:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_71_2914_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2932:142
    ._dfc_wire_104                          (_dup444__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:590:111
    ._dfc_wire_107                          (_MUL451__dfc_wire_107)
  );
  ADD_2x1 ADD452 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:598:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup449__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:595:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_163_2913_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2931:146
    ._dfc_wire_100                          (_ADD452__dfc_wire_100)
  );
  dup_1x2 dup453 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:599:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD428__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:574:130
    ._dfc_wire_68_105 (_dup453__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup453__dfc_wire_68_113)
  );
  dup_1x2 dup454 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:600:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB437__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:583:109
    ._dfc_wire_68_105 (_dup454__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup454__dfc_wire_68_113)
  );
  ADD_2x1 ADD455 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:601:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_72_2912_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2930:142
    .const_fix_32_0_1__0000000000000080_102 (_dup454__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:600:111
    ._dfc_wire_100                          (_ADD455__dfc_wire_100)
  );
  SUB_2x1 SUB456 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:602:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_72_2911_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2929:142
    ._dfc_wire_118    (_dup454__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:600:111
    ._dfc_wire_121    (_SUB456__dfc_wire_121)
  );
  dup_1x2 dup457 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:603:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB430__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:576:109
    ._dfc_wire_68_105 (_dup457__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup457__dfc_wire_68_113)
  );
  dup_1x2 dup458 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:604:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB439__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:585:109
    ._dfc_wire_68_105 (_dup458__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup458__dfc_wire_68_113)
  );
  ADD_2x1 ADD459 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:605:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_40_2910_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2928:142
    .const_fix_32_0_1__0000000000000080_102 (_dup458__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:604:111
    ._dfc_wire_100                          (_ADD459__dfc_wire_100)
  );
  SUB_2x1 SUB460 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:606:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_40_2909_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2927:142
    ._dfc_wire_118    (_dup458__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:604:111
    ._dfc_wire_121    (_SUB460__dfc_wire_121)
  );
  dup_1x2 dup461 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:607:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD442__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:588:130
    ._dfc_wire_68_105 (_dup461__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup461__dfc_wire_68_113)
  );
  dup_1x2 dup462 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:608:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD452__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:598:130
    ._dfc_wire_68_105 (_dup462__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup462__dfc_wire_68_113)
  );
  ADD_2x1 ADD463 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:609:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_45_2908_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2926:142
    .const_fix_32_0_1__0000000000000080_102 (_dup462__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:608:111
    ._dfc_wire_100                          (_ADD463__dfc_wire_100)
  );
  SUB_2x1 SUB464 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:610:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_45_2907_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2925:142
    ._dfc_wire_118    (_dup462__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:608:111
    ._dfc_wire_121    (_SUB464__dfc_wire_121)
  );
  dup_1x2 dup465 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:611:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB443__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:589:109
    ._dfc_wire_68_105 (_dup465__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup465__dfc_wire_68_113)
  );
  dup_1x2 dup466 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:612:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB450__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:596:109
    ._dfc_wire_68_105 (_dup466__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup466__dfc_wire_68_113)
  );
  ADD_2x1 ADD467 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:613:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup465__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:611:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_47_2906_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2924:142
    ._dfc_wire_100                          (_ADD467__dfc_wire_100)
  );
  SUB_2x1 SUB468 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:614:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup465__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:611:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_47_2905_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2923:142
    ._dfc_wire_121    (_SUB468__dfc_wire_121)
  );
  dup_1x2 dup469 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:615:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB456__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:602:109
    ._dfc_wire_68_105 (_dup469__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup469__dfc_wire_68_113)
  );
  dup_1x2 dup470 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:616:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB460__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:606:109
    ._dfc_wire_68_105 (_dup470__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup470__dfc_wire_68_113)
  );
  ADD_2x1 ADD471 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:617:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup469__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:615:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_103_2904_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2922:146
    ._dfc_wire_100                          (_ADD471__dfc_wire_100)
  );
  MUL_2x1 MUL472 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:618:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_504_2903_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2921:146
    ._dfc_wire_104                          (_ADD471__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:617:130
    ._dfc_wire_107                          (_MUL472__dfc_wire_107)
  );
  ADD_2x1 ADD473 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:619:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL472__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:618:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_605_2902_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2920:146
    ._dfc_wire_100                          (_ADD473__dfc_wire_100)
  );
  SHR8_1x1 SHR8474 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:620:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD473__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:619:130
    ._dfc_wire_216 (_SHR8474__dfc_wire_216)
  );
  SUB_2x1 SUB475 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:621:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup469__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:615:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_103_2901_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2919:146
    ._dfc_wire_121    (_SUB475__dfc_wire_121)
  );
  MUL_2x1 MUL476 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:622:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_473_2900_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2918:146
    ._dfc_wire_104                          (_SUB475__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:621:109
    ._dfc_wire_107                          (_MUL476__dfc_wire_107)
  );
  ADD_2x1 ADD477 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:623:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL476__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:622:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_561_2899_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2917:146
    ._dfc_wire_100                          (_ADD477__dfc_wire_100)
  );
  SHR8_1x1 SHR8478 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:624:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD477__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:623:130
    ._dfc_wire_216 (_SHR8478__dfc_wire_216)
  );
  dup_1x2 dup479 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:625:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD463__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:609:130
    ._dfc_wire_68_105 (_dup479__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup479__dfc_wire_68_113)
  );
  dup_1x2 dup480 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:626:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD455__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:601:130
    ._dfc_wire_68_105 (_dup480__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup480__dfc_wire_68_113)
  );
  ADD_2x1 ADD481 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:627:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_57_2898_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2916:142
    .const_fix_32_0_1__0000000000000080_102 (_dup480__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:626:111
    ._dfc_wire_100                          (_ADD481__dfc_wire_100)
  );
  SHR8_1x1 SHR8482 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:628:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD481__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:627:130
    ._dfc_wire_216 (_SHR8482__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST483 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:629:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8482__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:628:87
    ._dfc_wire_236 (_CAST483__dfc_wire_236)
  );
  dup_1x2 dup484 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:630:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD467__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:613:130
    ._dfc_wire_68_105 (_dup484__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup484__dfc_wire_68_113)
  );
  dup_1x2 dup485 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:631:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR8474__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:620:87
    ._dfc_wire_68_105 (_dup485__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup485__dfc_wire_68_113)
  );
  ADD_2x1 ADD486 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:632:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_272_2897_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2915:146
    .const_fix_32_0_1__0000000000000080_102 (_dup485__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:631:111
    ._dfc_wire_100                          (_ADD486__dfc_wire_100)
  );
  SHR8_1x1 SHR8487 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:633:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD486__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:632:130
    ._dfc_wire_216 (_SHR8487__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST488 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:634:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8487__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:633:87
    ._dfc_wire_236 (_CAST488__dfc_wire_236)
  );
  dup_1x2 dup489 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:635:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB468__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:614:109
    ._dfc_wire_68_105 (_dup489__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup489__dfc_wire_68_113)
  );
  dup_1x2 dup490 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:636:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR8478__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:624:87
    ._dfc_wire_68_105 (_dup490__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup490__dfc_wire_68_113)
  );
  ADD_2x1 ADD491 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:637:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_212_2896_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2914:146
    .const_fix_32_0_1__0000000000000080_102 (_dup490__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:636:111
    ._dfc_wire_100                          (_ADD491__dfc_wire_100)
  );
  SHR8_1x1 SHR8492 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:638:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD491__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:637:130
    ._dfc_wire_216 (_SHR8492__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST493 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:639:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8492__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:638:87
    ._dfc_wire_236 (_CAST493__dfc_wire_236)
  );
  dup_1x2 dup494 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:640:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB464__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:610:109
    ._dfc_wire_68_105 (_dup494__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup494__dfc_wire_68_113)
  );
  dup_1x2 dup495 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:641:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD459__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:605:130
    ._dfc_wire_68_105 (_dup495__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup495__dfc_wire_68_113)
  );
  ADD_2x1 ADD496 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:642:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup494__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:640:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_37_2895_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2913:142
    ._dfc_wire_100                          (_ADD496__dfc_wire_100)
  );
  SHR8_1x1 SHR8497 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:643:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD496__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:642:130
    ._dfc_wire_216 (_SHR8497__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST498 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:644:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8497__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:643:87
    ._dfc_wire_236 (_CAST498__dfc_wire_236)
  );
  SUB_2x1 SUB499 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:645:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup494__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:640:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_37_2894_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2912:142
    ._dfc_wire_121    (_SUB499__dfc_wire_121)
  );
  SHR8_1x1 SHR8500 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:646:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB499__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:645:109
    ._dfc_wire_216 (_SHR8500__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST501 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:647:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8500__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:646:87
    ._dfc_wire_236 (_CAST501__dfc_wire_236)
  );
  SUB_2x1 SUB502 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:648:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_212_2893_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2911:146
    ._dfc_wire_118    (_dup490__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:636:111
    ._dfc_wire_121    (_SUB502__dfc_wire_121)
  );
  SHR8_1x1 SHR8503 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:649:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB502__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:648:109
    ._dfc_wire_216 (_SHR8503__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST504 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:650:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8503__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:649:87
    ._dfc_wire_236 (_CAST504__dfc_wire_236)
  );
  SUB_2x1 SUB505 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:651:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_272_2892_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2910:146
    ._dfc_wire_118    (_dup485__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:631:111
    ._dfc_wire_121    (_SUB505__dfc_wire_121)
  );
  SHR8_1x1 SHR8506 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:652:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB505__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:651:109
    ._dfc_wire_216 (_SHR8506__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST507 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:653:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8506__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:652:87
    ._dfc_wire_236 (_CAST507__dfc_wire_236)
  );
  SUB_2x1 SUB508 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:654:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_57_2891_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2909:142
    ._dfc_wire_118    (_dup480__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:626:111
    ._dfc_wire_121    (_SUB508__dfc_wire_121)
  );
  SHR8_1x1 SHR8509 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:655:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB508__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:654:109
    ._dfc_wire_216 (_SHR8509__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST510 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:656:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8509__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:655:87
    ._dfc_wire_236 (_CAST510__dfc_wire_236)
  );
  CAST_1x1_16_32 CAST511 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:657:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_44__dfc_wire_45),
    ._dfc_wire_73 (_CAST511__dfc_wire_73)
  );
  SHL11_1x1 SHL11512 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:658:89
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_73 (_CAST511__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:657:84
    ._dfc_wire_75 (_SHL11512__dfc_wire_75)
  );
  CAST_1x1_16_32 CAST513 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:659:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_46__dfc_wire_45),
    ._dfc_wire_73 (_CAST513__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST514 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:660:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_42__dfc_wire_45),
    ._dfc_wire_73 (_CAST514__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST515 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:661:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_41__dfc_wire_45),
    ._dfc_wire_73 (_CAST515__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST516 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:662:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_47__dfc_wire_45),
    ._dfc_wire_73 (_CAST516__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST517 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:663:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_45__dfc_wire_45),
    ._dfc_wire_73 (_CAST517__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST518 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:664:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_43__dfc_wire_45),
    ._dfc_wire_73 (_CAST518__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST519 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:665:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_40__dfc_wire_45),
    ._dfc_wire_73 (_CAST519__dfc_wire_73)
  );
  SHL11_1x1 SHL11520 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:666:89
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_73 (_CAST519__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:665:84
    ._dfc_wire_75 (_SHL11520__dfc_wire_75)
  );
  ADD_2x1 ADD521 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:667:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_SHL11520__dfc_wire_75),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:666:89
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_132_2939_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2957:146
    ._dfc_wire_100                          (_ADD521__dfc_wire_100)
  );
  dup_1x2 dup522 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:668:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST515__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:661:84
    ._dfc_wire_68_105 (_dup522__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup522__dfc_wire_68_113)
  );
  dup_1x2 dup523 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:669:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST516__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:662:84
    ._dfc_wire_68_105 (_dup523__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup523__dfc_wire_68_113)
  );
  ADD_2x1 ADD524 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:670:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup522__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:668:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_10_2938_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2956:142
    ._dfc_wire_100                          (_ADD524__dfc_wire_100)
  );
  MUL_2x1 MUL525 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:671:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_162_2937_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2955:146
    ._dfc_wire_104                          (_ADD524__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:670:130
    ._dfc_wire_107                          (_MUL525__dfc_wire_107)
  );
  MUL_2x1 MUL526 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:672:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_75_2936_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2954:142
    ._dfc_wire_104                          (_dup522__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:668:111
    ._dfc_wire_107                          (_MUL526__dfc_wire_107)
  );
  dup_1x2 dup527 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:673:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL525__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:671:131
    ._dfc_wire_68_105 (_dup527__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup527__dfc_wire_68_113)
  );
  ADD_2x1 ADD528 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:674:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup527__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:673:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_57_2935_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2953:142
    ._dfc_wire_100                          (_ADD528__dfc_wire_100)
  );
  MUL_2x1 MUL529 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:675:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_109_2933_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2951:146
    ._dfc_wire_104                          (_dup523__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:669:111
    ._dfc_wire_107                          (_MUL529__dfc_wire_107)
  );
  SUB_2x1 SUB530 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:676:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup527__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:673:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_131_2890_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2908:146
    ._dfc_wire_121    (_SUB530__dfc_wire_121)
  );
  dup_1x2 dup531 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:677:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST517__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:663:84
    ._dfc_wire_68_105 (_dup531__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup531__dfc_wire_68_113)
  );
  dup_1x2 dup532 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:678:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST518__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:664:84
    ._dfc_wire_68_105 (_dup532__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup532__dfc_wire_68_113)
  );
  ADD_2x1 ADD533 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:679:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_70_2889_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2907:142
    .const_fix_32_0_1__0000000000000080_102 (_dup532__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:678:111
    ._dfc_wire_100                          (_ADD533__dfc_wire_100)
  );
  MUL_2x1 MUL534 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:680:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_145_2888_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2906:146
    ._dfc_wire_104                          (_ADD533__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:679:130
    ._dfc_wire_107                          (_MUL534__dfc_wire_107)
  );
  MUL_2x1 MUL535 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:681:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_10_2887_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2905:142
    ._dfc_wire_104                          (_dup531__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:677:111
    ._dfc_wire_107                          (_MUL535__dfc_wire_107)
  );
  dup_1x2 dup536 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:682:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL534__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:680:131
    ._dfc_wire_68_105 (_dup536__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup536__dfc_wire_68_113)
  );
  SUB_2x1 SUB537 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:683:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup536__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:682:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_103_2886_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2904:146
    ._dfc_wire_121    (_SUB537__dfc_wire_121)
  );
  MUL_2x1 MUL538 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:684:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_138_2885_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2903:146
    ._dfc_wire_104                          (_dup532__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:678:111
    ._dfc_wire_107                          (_MUL538__dfc_wire_107)
  );
  SUB_2x1 SUB539 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:685:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_3_2884_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2902:138
    ._dfc_wire_118    (_MUL538__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:684:131
    ._dfc_wire_121    (_SUB539__dfc_wire_121)
  );
  dup_1x2 dup540 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:686:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD521__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:667:130
    ._dfc_wire_68_105 (_dup540__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup540__dfc_wire_68_113)
  );
  dup_1x2 dup541 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:687:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHL11512__dfc_wire_75),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:658:89
    ._dfc_wire_68_105 (_dup541__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup541__dfc_wire_68_113)
  );
  ADD_2x1 ADD542 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:688:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup540__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:686:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_23_2883_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2901:142
    ._dfc_wire_100                          (_ADD542__dfc_wire_100)
  );
  SUB_2x1 SUB543 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:689:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup540__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:686:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_23_2882_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2900:142
    ._dfc_wire_121    (_SUB543__dfc_wire_121)
  );
  dup_1x2 dup544 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:690:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST514__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:660:84
    ._dfc_wire_68_105 (_dup544__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup544__dfc_wire_68_113)
  );
  dup_1x2 dup545 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:691:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST513__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:659:84
    ._dfc_wire_68_105 (_dup545__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup545__dfc_wire_68_113)
  );
  ADD_2x1 ADD546 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:692:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup544__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:690:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_2_2881_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2899:138
    ._dfc_wire_100                          (_ADD546__dfc_wire_100)
  );
  MUL_2x1 MUL547 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:693:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_177_2880_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2898:146
    ._dfc_wire_104                          (_ADD546__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:692:130
    ._dfc_wire_107                          (_MUL547__dfc_wire_107)
  );
  MUL_2x1 MUL548 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:694:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_64_2879_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2897:142
    ._dfc_wire_104                          (_dup545__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:691:111
    ._dfc_wire_107                          (_MUL548__dfc_wire_107)
  );
  dup_1x2 dup549 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:695:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL547__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:693:131
    ._dfc_wire_68_105 (_dup549__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup549__dfc_wire_68_113)
  );
  SUB_2x1 SUB550 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:696:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup549__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:695:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_110_2878_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2896:146
    ._dfc_wire_121    (_SUB550__dfc_wire_121)
  );
  MUL_2x1 MUL551 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:697:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_122_2877_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2895:146
    ._dfc_wire_104                          (_dup544__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:690:111
    ._dfc_wire_107                          (_MUL551__dfc_wire_107)
  );
  ADD_2x1 ADD552 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:698:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup549__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:695:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_95_2876_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2894:142
    ._dfc_wire_100                          (_ADD552__dfc_wire_100)
  );
  dup_1x2 dup553 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:699:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD528__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:674:130
    ._dfc_wire_68_105 (_dup553__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup553__dfc_wire_68_113)
  );
  dup_1x2 dup554 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:700:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB537__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:683:109
    ._dfc_wire_68_105 (_dup554__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup554__dfc_wire_68_113)
  );
  ADD_2x1 ADD555 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:701:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_1_2875_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2893:138
    .const_fix_32_0_1__0000000000000080_102 (_dup554__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:700:111
    ._dfc_wire_100                          (_ADD555__dfc_wire_100)
  );
  SUB_2x1 SUB556 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:702:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_1_2874_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2892:138
    ._dfc_wire_118    (_dup554__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:700:111
    ._dfc_wire_121    (_SUB556__dfc_wire_121)
  );
  dup_1x2 dup557 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:703:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB530__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:676:109
    ._dfc_wire_68_105 (_dup557__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup557__dfc_wire_68_113)
  );
  dup_1x2 dup558 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:704:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB539__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:685:109
    ._dfc_wire_68_105 (_dup558__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup558__dfc_wire_68_113)
  );
  ADD_2x1 ADD559 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:705:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup557__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:703:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_57_2873_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2891:142
    ._dfc_wire_100                          (_ADD559__dfc_wire_100)
  );
  SUB_2x1 SUB560 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:706:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup557__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:703:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_57_2872_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2890:142
    ._dfc_wire_121    (_SUB560__dfc_wire_121)
  );
  dup_1x2 dup561 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:707:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD542__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:688:130
    ._dfc_wire_68_105 (_dup561__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup561__dfc_wire_68_113)
  );
  dup_1x2 dup562 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:708:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD552__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:698:130
    ._dfc_wire_68_105 (_dup562__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup562__dfc_wire_68_113)
  );
  ADD_2x1 ADD563 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:709:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_118_2871_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2889:146
    .const_fix_32_0_1__0000000000000080_102 (_dup562__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:708:111
    ._dfc_wire_100                          (_ADD563__dfc_wire_100)
  );
  SUB_2x1 SUB564 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:710:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_118_2870_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2888:146
    ._dfc_wire_118    (_dup562__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:708:111
    ._dfc_wire_121    (_SUB564__dfc_wire_121)
  );
  dup_1x2 dup565 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:711:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB543__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:689:109
    ._dfc_wire_68_105 (_dup565__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup565__dfc_wire_68_113)
  );
  dup_1x2 dup566 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:712:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB550__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:696:109
    ._dfc_wire_68_105 (_dup566__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup566__dfc_wire_68_113)
  );
  ADD_2x1 ADD567 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:713:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_174_2869_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2887:146
    .const_fix_32_0_1__0000000000000080_102 (_dup566__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:712:111
    ._dfc_wire_100                          (_ADD567__dfc_wire_100)
  );
  SUB_2x1 SUB568 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:714:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_174_2868_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2886:146
    ._dfc_wire_118    (_dup566__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:712:111
    ._dfc_wire_121    (_SUB568__dfc_wire_121)
  );
  dup_1x2 dup569 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:715:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB556__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:702:109
    ._dfc_wire_68_105 (_dup569__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup569__dfc_wire_68_113)
  );
  dup_1x2 dup570 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:716:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB560__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:706:109
    ._dfc_wire_68_105 (_dup570__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup570__dfc_wire_68_113)
  );
  ADD_2x1 ADD571 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:717:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_94_2867_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2885:142
    .const_fix_32_0_1__0000000000000080_102 (_dup570__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:716:111
    ._dfc_wire_100                          (_ADD571__dfc_wire_100)
  );
  MUL_2x1 MUL572 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:718:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_497_2866_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2884:146
    ._dfc_wire_104                          (_ADD571__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:717:130
    ._dfc_wire_107                          (_MUL572__dfc_wire_107)
  );
  ADD_2x1 ADD573 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:719:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL572__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:718:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_610_2865_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2883:146
    ._dfc_wire_100                          (_ADD573__dfc_wire_100)
  );
  SHR8_1x1 SHR8574 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:720:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD573__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:719:130
    ._dfc_wire_216 (_SHR8574__dfc_wire_216)
  );
  SUB_2x1 SUB575 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:721:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_94_2864_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2882:142
    ._dfc_wire_118    (_dup570__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:716:111
    ._dfc_wire_121    (_SUB575__dfc_wire_121)
  );
  MUL_2x1 MUL576 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:722:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_516_2863_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2881:146
    ._dfc_wire_104                          (_SUB575__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:721:109
    ._dfc_wire_107                          (_MUL576__dfc_wire_107)
  );
  ADD_2x1 ADD577 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:723:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL576__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:722:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_670_2862_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2880:146
    ._dfc_wire_100                          (_ADD577__dfc_wire_100)
  );
  SHR8_1x1 SHR8578 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:724:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD577__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:723:130
    ._dfc_wire_216 (_SHR8578__dfc_wire_216)
  );
  dup_1x2 dup579 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:725:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD563__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:709:130
    ._dfc_wire_68_105 (_dup579__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup579__dfc_wire_68_113)
  );
  dup_1x2 dup580 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:726:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD555__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:701:130
    ._dfc_wire_68_105 (_dup580__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup580__dfc_wire_68_113)
  );
  ADD_2x1 ADD581 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:727:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_35_2861_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2879:142
    .const_fix_32_0_1__0000000000000080_102 (_dup580__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:726:111
    ._dfc_wire_100                          (_ADD581__dfc_wire_100)
  );
  SHR8_1x1 SHR8582 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:728:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD581__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:727:130
    ._dfc_wire_216 (_SHR8582__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST583 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:729:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8582__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:728:87
    ._dfc_wire_236 (_CAST583__dfc_wire_236)
  );
  dup_1x2 dup584 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:730:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD567__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:713:130
    ._dfc_wire_68_105 (_dup584__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup584__dfc_wire_68_113)
  );
  dup_1x2 dup585 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:731:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR8574__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:720:87
    ._dfc_wire_68_105 (_dup585__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup585__dfc_wire_68_113)
  );
  ADD_2x1 ADD586 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:732:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_134_2860_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2878:146
    .const_fix_32_0_1__0000000000000080_102 (_dup585__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:731:111
    ._dfc_wire_100                          (_ADD586__dfc_wire_100)
  );
  SHR8_1x1 SHR8587 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:733:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD586__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:732:130
    ._dfc_wire_216 (_SHR8587__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST588 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:734:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8587__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:733:87
    ._dfc_wire_236 (_CAST588__dfc_wire_236)
  );
  dup_1x2 dup589 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:735:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB568__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:714:109
    ._dfc_wire_68_105 (_dup589__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup589__dfc_wire_68_113)
  );
  dup_1x2 dup590 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:736:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR8578__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:724:87
    ._dfc_wire_68_105 (_dup590__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup590__dfc_wire_68_113)
  );
  ADD_2x1 ADD591 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:737:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_198_2859_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2877:146
    .const_fix_32_0_1__0000000000000080_102 (_dup590__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:736:111
    ._dfc_wire_100                          (_ADD591__dfc_wire_100)
  );
  SHR8_1x1 SHR8592 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:738:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD591__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:737:130
    ._dfc_wire_216 (_SHR8592__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST593 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:739:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8592__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:738:87
    ._dfc_wire_236 (_CAST593__dfc_wire_236)
  );
  dup_1x2 dup594 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:740:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB564__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:710:109
    ._dfc_wire_68_105 (_dup594__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup594__dfc_wire_68_113)
  );
  dup_1x2 dup595 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:741:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD559__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:705:130
    ._dfc_wire_68_105 (_dup595__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup595__dfc_wire_68_113)
  );
  ADD_2x1 ADD596 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:742:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup594__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:740:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_73_2858_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2876:142
    ._dfc_wire_100                          (_ADD596__dfc_wire_100)
  );
  SHR8_1x1 SHR8597 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:743:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD596__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:742:130
    ._dfc_wire_216 (_SHR8597__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST598 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:744:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8597__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:743:87
    ._dfc_wire_236 (_CAST598__dfc_wire_236)
  );
  SUB_2x1 SUB599 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:745:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup594__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:740:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_73_2857_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2875:142
    ._dfc_wire_121    (_SUB599__dfc_wire_121)
  );
  SHR8_1x1 SHR8600 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:746:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB599__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:745:109
    ._dfc_wire_216 (_SHR8600__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST601 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:747:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8600__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:746:87
    ._dfc_wire_236 (_CAST601__dfc_wire_236)
  );
  SUB_2x1 SUB602 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:748:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_198_2856_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2874:146
    ._dfc_wire_118    (_dup590__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:736:111
    ._dfc_wire_121    (_SUB602__dfc_wire_121)
  );
  SHR8_1x1 SHR8603 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:749:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB602__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:748:109
    ._dfc_wire_216 (_SHR8603__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST604 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:750:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8603__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:749:87
    ._dfc_wire_236 (_CAST604__dfc_wire_236)
  );
  SUB_2x1 SUB605 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:751:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_134_2855_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2873:146
    ._dfc_wire_118    (_dup585__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:731:111
    ._dfc_wire_121    (_SUB605__dfc_wire_121)
  );
  SHR8_1x1 SHR8606 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:752:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB605__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:751:109
    ._dfc_wire_216 (_SHR8606__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST607 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:753:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8606__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:752:87
    ._dfc_wire_236 (_CAST607__dfc_wire_236)
  );
  SUB_2x1 SUB608 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:754:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_35_2854_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2872:142
    ._dfc_wire_118    (_dup580__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:726:111
    ._dfc_wire_121    (_SUB608__dfc_wire_121)
  );
  SHR8_1x1 SHR8609 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:755:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB608__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:754:109
    ._dfc_wire_216 (_SHR8609__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST610 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:756:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8609__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:755:87
    ._dfc_wire_236 (_CAST610__dfc_wire_236)
  );
  CAST_1x1_16_32 CAST611 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:757:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_52__dfc_wire_45),
    ._dfc_wire_73 (_CAST611__dfc_wire_73)
  );
  SHL11_1x1 SHL11612 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:758:89
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_73 (_CAST611__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:757:84
    ._dfc_wire_75 (_SHL11612__dfc_wire_75)
  );
  CAST_1x1_16_32 CAST613 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:759:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_54__dfc_wire_45),
    ._dfc_wire_73 (_CAST613__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST614 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:760:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_50__dfc_wire_45),
    ._dfc_wire_73 (_CAST614__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST615 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:761:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_49__dfc_wire_45),
    ._dfc_wire_73 (_CAST615__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST616 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:762:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_55__dfc_wire_45),
    ._dfc_wire_73 (_CAST616__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST617 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:763:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_53__dfc_wire_45),
    ._dfc_wire_73 (_CAST617__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST618 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:764:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_51__dfc_wire_45),
    ._dfc_wire_73 (_CAST618__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST619 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:765:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_48__dfc_wire_45),
    ._dfc_wire_73 (_CAST619__dfc_wire_73)
  );
  SHL11_1x1 SHL11620 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:766:89
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_73 (_CAST619__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:765:84
    ._dfc_wire_75 (_SHL11620__dfc_wire_75)
  );
  ADD_2x1 ADD621 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:767:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_SHL11620__dfc_wire_75),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:766:89
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_113_2853_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2871:146
    ._dfc_wire_100                          (_ADD621__dfc_wire_100)
  );
  dup_1x2 dup622 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:768:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST615__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:761:84
    ._dfc_wire_68_105 (_dup622__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup622__dfc_wire_68_113)
  );
  dup_1x2 dup623 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:769:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST616__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:762:84
    ._dfc_wire_68_105 (_dup623__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup623__dfc_wire_68_113)
  );
  ADD_2x1 ADD624 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:770:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup622__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:768:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_73_2852_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2870:142
    ._dfc_wire_100                          (_ADD624__dfc_wire_100)
  );
  MUL_2x1 MUL625 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:771:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_202_2850_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2868:146
    ._dfc_wire_104                          (_ADD624__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:770:130
    ._dfc_wire_107                          (_MUL625__dfc_wire_107)
  );
  MUL_2x1 MUL626 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:772:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_175_2849_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2867:146
    ._dfc_wire_104                          (_dup622__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:768:111
    ._dfc_wire_107                          (_MUL626__dfc_wire_107)
  );
  dup_1x2 dup627 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:773:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL625__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:771:131
    ._dfc_wire_68_105 (_dup627__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup627__dfc_wire_68_113)
  );
  ADD_2x1 ADD628 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:774:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup627__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:773:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_24_2848_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2866:142
    ._dfc_wire_100                          (_ADD628__dfc_wire_100)
  );
  MUL_2x1 MUL629 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:775:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_146_2846_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2864:146
    ._dfc_wire_104                          (_dup623__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:769:111
    ._dfc_wire_107                          (_MUL629__dfc_wire_107)
  );
  SUB_2x1 SUB630 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:776:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup627__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:773:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_30_2844_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2862:142
    ._dfc_wire_121    (_SUB630__dfc_wire_121)
  );
  dup_1x2 dup631 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:777:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST617__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:763:84
    ._dfc_wire_68_105 (_dup631__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup631__dfc_wire_68_113)
  );
  dup_1x2 dup632 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:778:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST618__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:764:84
    ._dfc_wire_68_105 (_dup632__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup632__dfc_wire_68_113)
  );
  ADD_2x1 ADD633 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:779:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_29_2842_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2860:142
    .const_fix_32_0_1__0000000000000080_102 (_dup632__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:778:111
    ._dfc_wire_100                          (_ADD633__dfc_wire_100)
  );
  MUL_2x1 MUL634 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:780:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_164_2840_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2858:146
    ._dfc_wire_104                          (_ADD633__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:779:130
    ._dfc_wire_107                          (_MUL634__dfc_wire_107)
  );
  MUL_2x1 MUL635 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:781:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_40_2839_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2857:142
    ._dfc_wire_104                          (_dup631__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:777:111
    ._dfc_wire_107                          (_MUL635__dfc_wire_107)
  );
  dup_1x2 dup636 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:782:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL634__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:780:131
    ._dfc_wire_68_105 (_dup636__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup636__dfc_wire_68_113)
  );
  SUB_2x1 SUB637 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:783:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup636__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:782:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_61_2837_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2855:142
    ._dfc_wire_121    (_SUB637__dfc_wire_121)
  );
  MUL_2x1 MUL638 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:784:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_127_2835_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2853:146
    ._dfc_wire_104                          (_dup632__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:778:111
    ._dfc_wire_107                          (_MUL638__dfc_wire_107)
  );
  SUB_2x1 SUB639 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:785:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_11_2834_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2852:142
    ._dfc_wire_118    (_MUL638__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:784:131
    ._dfc_wire_121    (_SUB639__dfc_wire_121)
  );
  dup_1x2 dup640 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:786:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD621__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:767:130
    ._dfc_wire_68_105 (_dup640__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup640__dfc_wire_68_113)
  );
  dup_1x2 dup641 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:787:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHL11612__dfc_wire_75),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:758:89
    ._dfc_wire_68_105 (_dup641__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup641__dfc_wire_68_113)
  );
  ADD_2x1 ADD642 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:788:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup640__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:786:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_2_2831_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2849:138
    ._dfc_wire_100                          (_ADD642__dfc_wire_100)
  );
  SUB_2x1 SUB643 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:789:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup640__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:786:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_2_2830_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2848:138
    ._dfc_wire_121    (_SUB643__dfc_wire_121)
  );
  dup_1x2 dup644 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:790:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST614__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:760:84
    ._dfc_wire_68_105 (_dup644__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup644__dfc_wire_68_113)
  );
  dup_1x2 dup645 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:791:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST613__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:759:84
    ._dfc_wire_68_105 (_dup645__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup645__dfc_wire_68_113)
  );
  ADD_2x1 ADD646 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:792:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup644__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:790:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_129_2827_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2845:146
    ._dfc_wire_100                          (_ADD646__dfc_wire_100)
  );
  MUL_2x1 MUL647 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:793:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_229_2825_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2843:146
    ._dfc_wire_104                          (_ADD646__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:792:130
    ._dfc_wire_107                          (_MUL647__dfc_wire_107)
  );
  MUL_2x1 MUL648 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:794:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1_2824_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2842:138
    ._dfc_wire_104                          (_dup645__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:791:111
    ._dfc_wire_107                          (_MUL648__dfc_wire_107)
  );
  dup_1x2 dup649 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:795:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL647__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:793:131
    ._dfc_wire_68_105 (_dup649__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup649__dfc_wire_68_113)
  );
  SUB_2x1 SUB650 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:796:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup649__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:795:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_247_2821_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2839:146
    ._dfc_wire_121    (_SUB650__dfc_wire_121)
  );
  MUL_2x1 MUL651 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:797:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_186_2819_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2837:146
    ._dfc_wire_104                          (_dup644__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:790:111
    ._dfc_wire_107                          (_MUL651__dfc_wire_107)
  );
  ADD_2x1 ADD652 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:798:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup649__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:795:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_132_2818_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2836:146
    ._dfc_wire_100                          (_ADD652__dfc_wire_100)
  );
  dup_1x2 dup653 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:799:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD628__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:774:130
    ._dfc_wire_68_105 (_dup653__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup653__dfc_wire_68_113)
  );
  dup_1x2 dup654 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:800:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB637__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:783:109
    ._dfc_wire_68_105 (_dup654__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup654__dfc_wire_68_113)
  );
  ADD_2x1 ADD655 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:801:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_30_2816_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2834:142
    .const_fix_32_0_1__0000000000000080_102 (_dup654__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:800:111
    ._dfc_wire_100                          (_ADD655__dfc_wire_100)
  );
  SUB_2x1 SUB656 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:802:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_30_2815_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2833:142
    ._dfc_wire_118    (_dup654__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:800:111
    ._dfc_wire_121    (_SUB656__dfc_wire_121)
  );
  dup_1x2 dup657 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:803:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB630__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:776:109
    ._dfc_wire_68_105 (_dup657__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup657__dfc_wire_68_113)
  );
  dup_1x2 dup658 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:804:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB639__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:785:109
    ._dfc_wire_68_105 (_dup658__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup658__dfc_wire_68_113)
  );
  ADD_2x1 ADD659 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:805:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup657__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:803:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_7_2811_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2829:138
    ._dfc_wire_100                          (_ADD659__dfc_wire_100)
  );
  SUB_2x1 SUB660 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:806:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup657__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:803:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_7_2809_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2827:138
    ._dfc_wire_121    (_SUB660__dfc_wire_121)
  );
  dup_1x2 dup661 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:807:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD642__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:788:130
    ._dfc_wire_68_105 (_dup661__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup661__dfc_wire_68_113)
  );
  dup_1x2 dup662 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:808:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD652__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:798:130
    ._dfc_wire_68_105 (_dup662__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup662__dfc_wire_68_113)
  );
  ADD_2x1 ADD663 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:809:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_258_2806_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2824:146
    .const_fix_32_0_1__0000000000000080_102 (_dup662__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:808:111
    ._dfc_wire_100                          (_ADD663__dfc_wire_100)
  );
  SUB_2x1 SUB664 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:810:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_258_2805_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2823:146
    ._dfc_wire_118    (_dup662__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:808:111
    ._dfc_wire_121    (_SUB664__dfc_wire_121)
  );
  dup_1x2 dup665 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:811:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB643__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:789:109
    ._dfc_wire_68_105 (_dup665__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup665__dfc_wire_68_113)
  );
  dup_1x2 dup666 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:812:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB650__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:796:109
    ._dfc_wire_68_105 (_dup666__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup666__dfc_wire_68_113)
  );
  ADD_2x1 ADD667 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:813:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_177_2803_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2821:146
    .const_fix_32_0_1__0000000000000080_102 (_dup666__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:812:111
    ._dfc_wire_100                          (_ADD667__dfc_wire_100)
  );
  SUB_2x1 SUB668 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:814:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_177_2801_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2819:146
    ._dfc_wire_118    (_dup666__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:812:111
    ._dfc_wire_121    (_SUB668__dfc_wire_121)
  );
  dup_1x2 dup669 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:815:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB656__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:802:109
    ._dfc_wire_68_105 (_dup669__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup669__dfc_wire_68_113)
  );
  dup_1x2 dup670 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:816:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB660__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:806:109
    ._dfc_wire_68_105 (_dup670__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup670__dfc_wire_68_113)
  );
  ADD_2x1 ADD671 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:817:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup669__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:815:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_98_2795_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2813:142
    ._dfc_wire_100                          (_ADD671__dfc_wire_100)
  );
  MUL_2x1 MUL672 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:818:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_417_2794_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2812:146
    ._dfc_wire_104                          (_ADD671__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:817:130
    ._dfc_wire_107                          (_MUL672__dfc_wire_107)
  );
  ADD_2x1 ADD673 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:819:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL672__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:818:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_584_2793_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2811:146
    ._dfc_wire_100                          (_ADD673__dfc_wire_100)
  );
  SHR8_1x1 SHR8674 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:820:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD673__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:819:130
    ._dfc_wire_216 (_SHR8674__dfc_wire_216)
  );
  SUB_2x1 SUB675 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:821:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup669__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:815:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_98_2791_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2809:142
    ._dfc_wire_121    (_SUB675__dfc_wire_121)
  );
  MUL_2x1 MUL676 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:822:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_442_2790_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2808:146
    ._dfc_wire_104                          (_SUB675__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:821:109
    ._dfc_wire_107                          (_MUL676__dfc_wire_107)
  );
  ADD_2x1 ADD677 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:823:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL676__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:822:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_537_2789_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2807:146
    ._dfc_wire_100                          (_ADD677__dfc_wire_100)
  );
  SHR8_1x1 SHR8678 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:824:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD677__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:823:130
    ._dfc_wire_216 (_SHR8678__dfc_wire_216)
  );
  dup_1x2 dup679 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:825:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD663__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:809:130
    ._dfc_wire_68_105 (_dup679__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup679__dfc_wire_68_113)
  );
  dup_1x2 dup680 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:826:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD655__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:801:130
    ._dfc_wire_68_105 (_dup680__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup680__dfc_wire_68_113)
  );
  ADD_2x1 ADD681 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:827:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup679__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:825:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_90_2782_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2800:142
    ._dfc_wire_100                          (_ADD681__dfc_wire_100)
  );
  SHR8_1x1 SHR8682 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:828:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD681__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:827:130
    ._dfc_wire_216 (_SHR8682__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST683 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:829:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8682__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:828:87
    ._dfc_wire_236 (_CAST683__dfc_wire_236)
  );
  dup_1x2 dup684 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:830:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD667__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:813:130
    ._dfc_wire_68_105 (_dup684__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup684__dfc_wire_68_113)
  );
  dup_1x2 dup685 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:831:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR8674__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:820:87
    ._dfc_wire_68_105 (_dup685__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup685__dfc_wire_68_113)
  );
  ADD_2x1 ADD686 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:832:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_65_2780_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2798:142
    .const_fix_32_0_1__0000000000000080_102 (_dup685__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:831:111
    ._dfc_wire_100                          (_ADD686__dfc_wire_100)
  );
  SHR8_1x1 SHR8687 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:833:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD686__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:832:130
    ._dfc_wire_216 (_SHR8687__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST688 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:834:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8687__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:833:87
    ._dfc_wire_236 (_CAST688__dfc_wire_236)
  );
  dup_1x2 dup689 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:835:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB668__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:814:109
    ._dfc_wire_68_105 (_dup689__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup689__dfc_wire_68_113)
  );
  dup_1x2 dup690 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:836:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR8678__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:824:87
    ._dfc_wire_68_105 (_dup690__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup690__dfc_wire_68_113)
  );
  ADD_2x1 ADD691 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:837:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_249_2773_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2791:146
    .const_fix_32_0_1__0000000000000080_102 (_dup690__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:836:111
    ._dfc_wire_100                          (_ADD691__dfc_wire_100)
  );
  SHR8_1x1 SHR8692 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:838:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD691__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:837:130
    ._dfc_wire_216 (_SHR8692__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST693 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:839:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8692__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:838:87
    ._dfc_wire_236 (_CAST693__dfc_wire_236)
  );
  dup_1x2 dup694 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:840:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB664__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:810:109
    ._dfc_wire_68_105 (_dup694__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup694__dfc_wire_68_113)
  );
  dup_1x2 dup695 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:841:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD659__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:805:130
    ._dfc_wire_68_105 (_dup695__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup695__dfc_wire_68_113)
  );
  ADD_2x1 ADD696 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:842:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup694__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:840:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_108_2770_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2788:146
    ._dfc_wire_100                          (_ADD696__dfc_wire_100)
  );
  SHR8_1x1 SHR8697 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:843:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD696__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:842:130
    ._dfc_wire_216 (_SHR8697__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST698 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:844:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8697__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:843:87
    ._dfc_wire_236 (_CAST698__dfc_wire_236)
  );
  SUB_2x1 SUB699 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:845:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup694__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:840:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_108_2764_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2782:146
    ._dfc_wire_121    (_SUB699__dfc_wire_121)
  );
  SHR8_1x1 SHR8700 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:846:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB699__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:845:109
    ._dfc_wire_216 (_SHR8700__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST701 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:847:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8700__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:846:87
    ._dfc_wire_236 (_CAST701__dfc_wire_236)
  );
  SUB_2x1 SUB702 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:848:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_249_2762_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2780:146
    ._dfc_wire_118    (_dup690__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:836:111
    ._dfc_wire_121    (_SUB702__dfc_wire_121)
  );
  SHR8_1x1 SHR8703 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:849:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB702__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:848:109
    ._dfc_wire_216 (_SHR8703__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST704 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:850:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8703__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:849:87
    ._dfc_wire_236 (_CAST704__dfc_wire_236)
  );
  SUB_2x1 SUB705 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:851:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_65_2758_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2776:142
    ._dfc_wire_118    (_dup685__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:831:111
    ._dfc_wire_121    (_SUB705__dfc_wire_121)
  );
  SHR8_1x1 SHR8706 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:852:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB705__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:851:109
    ._dfc_wire_216 (_SHR8706__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST707 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:853:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8706__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:852:87
    ._dfc_wire_236 (_CAST707__dfc_wire_236)
  );
  SUB_2x1 SUB708 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:854:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup679__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:825:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_90_2754_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2772:142
    ._dfc_wire_121    (_SUB708__dfc_wire_121)
  );
  SHR8_1x1 SHR8709 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:855:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB708__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:854:109
    ._dfc_wire_216 (_SHR8709__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST710 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:856:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8709__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:855:87
    ._dfc_wire_236 (_CAST710__dfc_wire_236)
  );
  CAST_1x1_16_32 CAST711 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:857:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_60__dfc_wire_45),
    ._dfc_wire_73 (_CAST711__dfc_wire_73)
  );
  SHL11_1x1 SHL11712 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:858:89
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_73 (_CAST711__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:857:84
    ._dfc_wire_75 (_SHL11712__dfc_wire_75)
  );
  CAST_1x1_16_32 CAST713 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:859:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_62__dfc_wire_45),
    ._dfc_wire_73 (_CAST713__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST714 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:860:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_58__dfc_wire_45),
    ._dfc_wire_73 (_CAST714__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST715 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:861:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_57__dfc_wire_45),
    ._dfc_wire_73 (_CAST715__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST716 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:862:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_63__dfc_wire_45),
    ._dfc_wire_73 (_CAST716__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST717 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:863:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_61__dfc_wire_45),
    ._dfc_wire_73 (_CAST717__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST718 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:864:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_59__dfc_wire_45),
    ._dfc_wire_73 (_CAST718__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST719 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:865:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (source__dfc_wire_56__dfc_wire_45),
    ._dfc_wire_73 (_CAST719__dfc_wire_73)
  );
  SHL11_1x1 SHL11720 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:866:89
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_73 (_CAST719__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:865:84
    ._dfc_wire_75 (_SHL11720__dfc_wire_75)
  );
  ADD_2x1 ADD721 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:867:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_SHL11720__dfc_wire_75),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:866:89
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_134_2742_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2760:146
    ._dfc_wire_100                          (_ADD721__dfc_wire_100)
  );
  dup_1x2 dup722 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:868:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST715__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:861:84
    ._dfc_wire_68_105 (_dup722__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup722__dfc_wire_68_113)
  );
  dup_1x2 dup723 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:869:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST716__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:862:84
    ._dfc_wire_68_105 (_dup723__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup723__dfc_wire_68_113)
  );
  ADD_2x1 ADD724 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:870:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_13_2738_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2756:142
    .const_fix_32_0_1__0000000000000080_102 (_dup723__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:869:111
    ._dfc_wire_100                          (_ADD724__dfc_wire_100)
  );
  MUL_2x1 MUL725 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:871:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_75_2737_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2755:142
    ._dfc_wire_104                          (_ADD724__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:870:130
    ._dfc_wire_107                          (_MUL725__dfc_wire_107)
  );
  MUL_2x1 MUL726 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:872:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_dup17_const_fix_32_0_1__0000000000000235_1725),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
    ._dfc_wire_104                          (_delay_fixed_32_0_1_4_2736_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2754:138
    ._dfc_wire_107                          (_MUL726__dfc_wire_107)
  );
  dup_1x2 dup727 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:873:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL725__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:871:131
    ._dfc_wire_68_105 (_dup727__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup727__dfc_wire_68_113)
  );
  ADD_2x1 ADD728 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:874:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup727__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:873:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_88_2735_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2753:142
    ._dfc_wire_100                          (_ADD728__dfc_wire_100)
  );
  MUL_2x1 MUL729 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:875:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_53_2734_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2752:142
    ._dfc_wire_104                          (_dup723__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:869:111
    ._dfc_wire_107                          (_MUL729__dfc_wire_107)
  );
  SUB_2x1 SUB730 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:876:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup727__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:873:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_122_2733_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2751:146
    ._dfc_wire_121    (_SUB730__dfc_wire_121)
  );
  dup_1x2 dup731 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:877:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST717__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:863:84
    ._dfc_wire_68_105 (_dup731__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup731__dfc_wire_68_113)
  );
  dup_1x2 dup732 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:878:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST718__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:864:84
    ._dfc_wire_68_105 (_dup732__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup732__dfc_wire_68_113)
  );
  ADD_2x1 ADD733 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:879:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_82_2732_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2750:142
    .const_fix_32_0_1__0000000000000080_102 (_dup732__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:878:111
    ._dfc_wire_100                          (_ADD733__dfc_wire_100)
  );
  MUL_2x1 MUL734 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:880:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_124_2731_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2749:146
    ._dfc_wire_104                          (_ADD733__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:879:130
    ._dfc_wire_107                          (_MUL734__dfc_wire_107)
  );
  MUL_2x1 MUL735 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:881:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_dup29_const_fix_32_0_1__0000000000000235_1725),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
    ._dfc_wire_104                          (_delay_fixed_32_0_1_21_2729_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2747:142
    ._dfc_wire_107                          (_MUL735__dfc_wire_107)
  );
  dup_1x2 dup736 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:882:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL734__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:880:131
    ._dfc_wire_68_105 (_dup736__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup736__dfc_wire_68_113)
  );
  SUB_2x1 SUB737 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:883:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup736__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:882:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_131_2728_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2746:146
    ._dfc_wire_121    (_SUB737__dfc_wire_121)
  );
  MUL_2x1 MUL738 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:884:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_119_2726_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2744:146
    ._dfc_wire_104                          (_dup732__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:878:111
    ._dfc_wire_107                          (_MUL738__dfc_wire_107)
  );
  SUB_2x1 SUB739 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:885:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup736__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:882:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_17_2724_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2742:142
    ._dfc_wire_121    (_SUB739__dfc_wire_121)
  );
  dup_1x2 dup740 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:886:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD721__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:867:130
    ._dfc_wire_68_105 (_dup740__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup740__dfc_wire_68_113)
  );
  dup_1x2 dup741 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:887:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHL11712__dfc_wire_75),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:858:89
    ._dfc_wire_68_105 (_dup741__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup741__dfc_wire_68_113)
  );
  ADD_2x1 ADD742 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:888:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup740__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:886:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_3_2720_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2738:138
    ._dfc_wire_100                          (_ADD742__dfc_wire_100)
  );
  SUB_2x1 SUB743 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:889:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup740__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:886:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_3_2716_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2734:138
    ._dfc_wire_121    (_SUB743__dfc_wire_121)
  );
  dup_1x2 dup744 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:890:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST714__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:860:84
    ._dfc_wire_68_105 (_dup744__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup744__dfc_wire_68_113)
  );
  dup_1x2 dup745 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:891:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST713__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:859:84
    ._dfc_wire_68_105 (_dup745__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup745__dfc_wire_68_113)
  );
  ADD_2x1 ADD746 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:892:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_80_2710_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2728:142
    .const_fix_32_0_1__0000000000000080_102 (_dup745__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:891:111
    ._dfc_wire_100                          (_ADD746__dfc_wire_100)
  );
  MUL_2x1 MUL747 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:893:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_155_2709_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2727:146
    ._dfc_wire_104                          (_ADD746__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:892:130
    ._dfc_wire_107                          (_MUL747__dfc_wire_107)
  );
  MUL_2x1 MUL748 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:894:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_98_2708_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2726:142
    ._dfc_wire_104                          (_dup745__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:891:111
    ._dfc_wire_107                          (_MUL748__dfc_wire_107)
  );
  dup_1x2 dup749 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:895:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_MUL747__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:893:131
    ._dfc_wire_68_105 (_dup749__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup749__dfc_wire_68_113)
  );
  SUB_2x1 SUB750 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:896:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup749__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:895:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_141_2705_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2723:146
    ._dfc_wire_121    (_SUB750__dfc_wire_121)
  );
  MUL_2x1 MUL751 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:897:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_74_2703_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2721:142
    ._dfc_wire_104                          (_dup744__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:890:111
    ._dfc_wire_107                          (_MUL751__dfc_wire_107)
  );
  ADD_2x1 ADD752 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:898:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup749__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:895:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_198_2701_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2719:146
    ._dfc_wire_100                          (_ADD752__dfc_wire_100)
  );
  dup_1x2 dup753 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:899:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD728__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:874:130
    ._dfc_wire_68_105 (_dup753__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup753__dfc_wire_68_113)
  );
  dup_1x2 dup754 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:900:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB737__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:883:109
    ._dfc_wire_68_105 (_dup754__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup754__dfc_wire_68_113)
  );
  ADD_2x1 ADD755 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:901:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup753__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:899:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_135_2694_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2712:146
    ._dfc_wire_100                          (_ADD755__dfc_wire_100)
  );
  SUB_2x1 SUB756 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:902:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup753__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:899:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_135_2691_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2709:146
    ._dfc_wire_121    (_SUB756__dfc_wire_121)
  );
  dup_1x2 dup757 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:903:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB730__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:876:109
    ._dfc_wire_68_105 (_dup757__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup757__dfc_wire_68_113)
  );
  dup_1x2 dup758 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:904:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB739__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:885:109
    ._dfc_wire_68_105 (_dup758__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup758__dfc_wire_68_113)
  );
  ADD_2x1 ADD759 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:905:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_1_2688_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2706:138
    .const_fix_32_0_1__0000000000000080_102 (_dup758__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:904:111
    ._dfc_wire_100                          (_ADD759__dfc_wire_100)
  );
  SUB_2x1 SUB760 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:906:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_1_2686_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2704:138
    ._dfc_wire_118    (_dup758__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:904:111
    ._dfc_wire_121    (_SUB760__dfc_wire_121)
  );
  dup_1x2 dup761 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:907:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD742__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:888:130
    ._dfc_wire_68_105 (_dup761__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup761__dfc_wire_68_113)
  );
  dup_1x2 dup762 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:908:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD752__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:898:130
    ._dfc_wire_68_105 (_dup762__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup762__dfc_wire_68_113)
  );
  ADD_2x1 ADD763 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:909:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_55_2682_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2700:142
    .const_fix_32_0_1__0000000000000080_102 (_dup762__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:908:111
    ._dfc_wire_100                          (_ADD763__dfc_wire_100)
  );
  SUB_2x1 SUB764 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:910:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_55_2679_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2697:142
    ._dfc_wire_118    (_dup762__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:908:111
    ._dfc_wire_121    (_SUB764__dfc_wire_121)
  );
  dup_1x2 dup765 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:911:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB743__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:889:109
    ._dfc_wire_68_105 (_dup765__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup765__dfc_wire_68_113)
  );
  dup_1x2 dup766 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:912:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB750__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:896:109
    ._dfc_wire_68_105 (_dup766__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup766__dfc_wire_68_113)
  );
  ADD_2x1 ADD767 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:913:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_50_2673_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2691:142
    .const_fix_32_0_1__0000000000000080_102 (_dup766__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:912:111
    ._dfc_wire_100                          (_ADD767__dfc_wire_100)
  );
  SUB_2x1 SUB768 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:914:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_50_2671_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2689:142
    ._dfc_wire_118    (_dup766__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:912:111
    ._dfc_wire_121    (_SUB768__dfc_wire_121)
  );
  dup_1x2 dup769 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:915:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB756__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:902:109
    ._dfc_wire_68_105 (_dup769__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup769__dfc_wire_68_113)
  );
  dup_1x2 dup770 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:916:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB760__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:906:109
    ._dfc_wire_68_105 (_dup770__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup770__dfc_wire_68_113)
  );
  ADD_2x1 ADD771 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:917:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_12_2667_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2685:142
    .const_fix_32_0_1__0000000000000080_102 (_dup770__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:916:111
    ._dfc_wire_100                          (_ADD771__dfc_wire_100)
  );
  MUL_2x1 MUL772 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:918:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_472_2666_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2684:146
    ._dfc_wire_104                          (_ADD771__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:917:130
    ._dfc_wire_107                          (_MUL772__dfc_wire_107)
  );
  ADD_2x1 ADD773 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:919:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL772__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:918:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_552_2663_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2681:146
    ._dfc_wire_100                          (_ADD773__dfc_wire_100)
  );
  SHR8_1x1 SHR8774 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:920:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD773__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:919:130
    ._dfc_wire_216 (_SHR8774__dfc_wire_216)
  );
  SUB_2x1 SUB775 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:921:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_12_2658_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2676:142
    ._dfc_wire_118    (_dup770__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:916:111
    ._dfc_wire_121    (_SUB775__dfc_wire_121)
  );
  MUL_2x1 MUL776 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:922:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_473_2655_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2673:146
    ._dfc_wire_104                          (_SUB775__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:921:109
    ._dfc_wire_107                          (_MUL776__dfc_wire_107)
  );
  ADD_2x1 ADD777 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:923:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL776__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:922:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_622_2654_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2672:146
    ._dfc_wire_100                          (_ADD777__dfc_wire_100)
  );
  SHR8_1x1 SHR8778 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:924:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD777__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:923:130
    ._dfc_wire_216 (_SHR8778__dfc_wire_216)
  );
  dup_1x2 dup779 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:925:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD763__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:909:130
    ._dfc_wire_68_105 (_dup779__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup779__dfc_wire_68_113)
  );
  dup_1x2 dup780 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:926:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD755__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:901:130
    ._dfc_wire_68_105 (_dup780__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup780__dfc_wire_68_113)
  );
  ADD_2x1 ADD781 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:927:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_85_2649_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2667:142
    .const_fix_32_0_1__0000000000000080_102 (_dup780__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:926:111
    ._dfc_wire_100                          (_ADD781__dfc_wire_100)
  );
  SHR8_1x1 SHR8782 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:928:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD781__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:927:130
    ._dfc_wire_216 (_SHR8782__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST783 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:929:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8782__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:928:87
    ._dfc_wire_236 (_CAST783__dfc_wire_236)
  );
  dup_1x2 dup784 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:930:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD767__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:913:130
    ._dfc_wire_68_105 (_dup784__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup784__dfc_wire_68_113)
  );
  dup_1x2 dup785 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:931:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR8774__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:920:87
    ._dfc_wire_68_105 (_dup785__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup785__dfc_wire_68_113)
  );
  ADD_2x1 ADD786 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:932:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_149_2643_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2661:146
    .const_fix_32_0_1__0000000000000080_102 (_dup785__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:931:111
    ._dfc_wire_100                          (_ADD786__dfc_wire_100)
  );
  SHR8_1x1 SHR8787 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:933:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD786__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:932:130
    ._dfc_wire_216 (_SHR8787__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST788 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:934:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8787__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:933:87
    ._dfc_wire_236 (_CAST788__dfc_wire_236)
  );
  dup_1x2 dup789 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:935:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB768__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:914:109
    ._dfc_wire_68_105 (_dup789__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup789__dfc_wire_68_113)
  );
  dup_1x2 dup790 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:936:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR8778__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:924:87
    ._dfc_wire_68_105 (_dup790__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup790__dfc_wire_68_113)
  );
  ADD_2x1 ADD791 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:937:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_151_2639_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2657:146
    .const_fix_32_0_1__0000000000000080_102 (_dup790__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:936:111
    ._dfc_wire_100                          (_ADD791__dfc_wire_100)
  );
  SHR8_1x1 SHR8792 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:938:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD791__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:937:130
    ._dfc_wire_216 (_SHR8792__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST793 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:939:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8792__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:938:87
    ._dfc_wire_236 (_CAST793__dfc_wire_236)
  );
  dup_1x2 dup794 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:940:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB764__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:910:109
    ._dfc_wire_68_105 (_dup794__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup794__dfc_wire_68_113)
  );
  dup_1x2 dup795 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:941:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD759__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:905:130
    ._dfc_wire_68_105 (_dup795__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup795__dfc_wire_68_113)
  );
  ADD_2x1 ADD796 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:942:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup794__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:940:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_22_2635_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2653:142
    ._dfc_wire_100                          (_ADD796__dfc_wire_100)
  );
  SHR8_1x1 SHR8797 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:943:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD796__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:942:130
    ._dfc_wire_216 (_SHR8797__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST798 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:944:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8797__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:943:87
    ._dfc_wire_236 (_CAST798__dfc_wire_236)
  );
  SUB_2x1 SUB799 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:945:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup794__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:940:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_22_2632_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2650:142
    ._dfc_wire_121    (_SUB799__dfc_wire_121)
  );
  SHR8_1x1 SHR8800 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:946:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB799__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:945:109
    ._dfc_wire_216 (_SHR8800__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST801 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:947:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8800__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:946:87
    ._dfc_wire_236 (_CAST801__dfc_wire_236)
  );
  SUB_2x1 SUB802 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:948:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_151_2627_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2645:146
    ._dfc_wire_118    (_dup790__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:936:111
    ._dfc_wire_121    (_SUB802__dfc_wire_121)
  );
  SHR8_1x1 SHR8803 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:949:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB802__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:948:109
    ._dfc_wire_216 (_SHR8803__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST804 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:950:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8803__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:949:87
    ._dfc_wire_236 (_CAST804__dfc_wire_236)
  );
  SUB_2x1 SUB805 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:951:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_149_2624_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2642:146
    ._dfc_wire_118    (_dup785__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:931:111
    ._dfc_wire_121    (_SUB805__dfc_wire_121)
  );
  SHR8_1x1 SHR8806 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:952:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB805__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:951:109
    ._dfc_wire_216 (_SHR8806__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST807 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:953:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8806__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:952:87
    ._dfc_wire_236 (_CAST807__dfc_wire_236)
  );
  SUB_2x1 SUB808 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:954:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_85_2617_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2635:142
    ._dfc_wire_118    (_dup780__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:926:111
    ._dfc_wire_121    (_SUB808__dfc_wire_121)
  );
  SHR8_1x1 SHR8809 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:955:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_SUB808__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:954:109
    ._dfc_wire_216 (_SHR8809__dfc_wire_216)
  );
  CAST_1x1_32_16 CAST810 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:956:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_SHR8809__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:955:87
    ._dfc_wire_236 (_CAST810__dfc_wire_236)
  );
  CAST_1x1_16_32 CAST811 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:957:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST483__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:629:87
    ._dfc_wire_73 (_CAST811__dfc_wire_73)
  );
  SHL8_1x1 SHL8812 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:958:89
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1921 (_CAST811__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:957:84
    ._dfc_wire_1923 (_SHL8812__dfc_wire_1923)
  );
  CAST_1x1_16_32 CAST813 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:959:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST683__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:829:87
    ._dfc_wire_73 (_CAST813__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST814 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:960:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST283__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:429:87
    ._dfc_wire_73 (_CAST814__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST815 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:961:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST183__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:329:87
    ._dfc_wire_73 (_CAST815__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST816 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:962:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST783__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:929:87
    ._dfc_wire_73 (_CAST816__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST817 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:963:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST583__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:729:87
    ._dfc_wire_73 (_CAST817__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST818 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:964:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST383__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:529:87
    ._dfc_wire_73 (_CAST818__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST819 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:965:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST83__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:229:83
    ._dfc_wire_73 (_CAST819__dfc_wire_73)
  );
  SHL8_1x1 SHL8820 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:966:89
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1921 (_CAST819__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:965:84
    ._dfc_wire_1923 (_SHL8820__dfc_wire_1923)
  );
  dup_1x8 dup821 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:967:473
    .clock                                   (clock),
    .reset                                   (reset),
    .const_fix_32_0_1__0000000000002000      (_const2045_const_fix_32_0_1__0000000000002000),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2153:90
    .const_fix_32_0_1__0000000000002000_1950 (_dup821_const_fix_32_0_1__0000000000002000_1950),
    .const_fix_32_0_1__0000000000002000_2314 (_dup821_const_fix_32_0_1__0000000000002000_2314),
    .const_fix_32_0_1__0000000000002000_2678 (_dup821_const_fix_32_0_1__0000000000002000_2678),
    .const_fix_32_0_1__0000000000002000_3042 (_dup821_const_fix_32_0_1__0000000000002000_3042),
    .const_fix_32_0_1__0000000000002000_3406 (_dup821_const_fix_32_0_1__0000000000002000_3406),
    .const_fix_32_0_1__0000000000002000_3770 (_dup821_const_fix_32_0_1__0000000000002000_3770),
    .const_fix_32_0_1__0000000000002000_4134 (_dup821_const_fix_32_0_1__0000000000002000_4134),
    .const_fix_32_0_1__0000000000002000_4498 (_dup821_const_fix_32_0_1__0000000000002000_4498)
  );
  ADD_2x1 ADD822 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:968:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_SHL8820__dfc_wire_1923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:966:89
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_825_2595_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2613:146
    ._dfc_wire_100                          (_ADD822__dfc_wire_100)
  );
  dup_1x2 dup823 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:969:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST815__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:961:84
    ._dfc_wire_68_105 (_dup823__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup823__dfc_wire_68_113)
  );
  dup_1x2 dup824 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:970:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST816__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:962:84
    ._dfc_wire_68_105 (_dup824__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup824__dfc_wire_68_113)
  );
  ADD_2x1 ADD825 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:971:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup823__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:969:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_41_2589_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2607:142
    ._dfc_wire_100                          (_ADD825__dfc_wire_100)
  );
  MUL_2x1 MUL826 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:972:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_744_2586_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2604:146
    ._dfc_wire_104                          (_ADD825__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:971:130
    ._dfc_wire_107                          (_MUL826__dfc_wire_107)
  );
  dup_1x24 dup827 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .clock                                   (clock),
    .reset                                   (reset),
    .const_fix_32_0_1__0000000000000004      (_const2144_const_fix_32_0_1__0000000000000004),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2165:90
    .const_fix_32_0_1__0000000000000004_1960 (_dup827_const_fix_32_0_1__0000000000000004_1960),
    .const_fix_32_0_1__0000000000000004_1988 (_dup827_const_fix_32_0_1__0000000000000004_1988),
    .const_fix_32_0_1__0000000000000004_2024 (_dup827_const_fix_32_0_1__0000000000000004_2024),
    .const_fix_32_0_1__0000000000000004_2324 (_dup827_const_fix_32_0_1__0000000000000004_2324),
    .const_fix_32_0_1__0000000000000004_2352 (_dup827_const_fix_32_0_1__0000000000000004_2352),
    .const_fix_32_0_1__0000000000000004_2388 (_dup827_const_fix_32_0_1__0000000000000004_2388),
    .const_fix_32_0_1__0000000000000004_2688 (_dup827_const_fix_32_0_1__0000000000000004_2688),
    .const_fix_32_0_1__0000000000000004_2716 (_dup827_const_fix_32_0_1__0000000000000004_2716),
    .const_fix_32_0_1__0000000000000004_2752 (_dup827_const_fix_32_0_1__0000000000000004_2752),
    .const_fix_32_0_1__0000000000000004_3052 (_dup827_const_fix_32_0_1__0000000000000004_3052),
    .const_fix_32_0_1__0000000000000004_3080 (_dup827_const_fix_32_0_1__0000000000000004_3080),
    .const_fix_32_0_1__0000000000000004_3116 (_dup827_const_fix_32_0_1__0000000000000004_3116),
    .const_fix_32_0_1__0000000000000004_3416 (_dup827_const_fix_32_0_1__0000000000000004_3416),
    .const_fix_32_0_1__0000000000000004_3444 (_dup827_const_fix_32_0_1__0000000000000004_3444),
    .const_fix_32_0_1__0000000000000004_3480 (_dup827_const_fix_32_0_1__0000000000000004_3480),
    .const_fix_32_0_1__0000000000000004_3780 (_dup827_const_fix_32_0_1__0000000000000004_3780),
    .const_fix_32_0_1__0000000000000004_3808 (_dup827_const_fix_32_0_1__0000000000000004_3808),
    .const_fix_32_0_1__0000000000000004_3844 (_dup827_const_fix_32_0_1__0000000000000004_3844),
    .const_fix_32_0_1__0000000000000004_4144 (_dup827_const_fix_32_0_1__0000000000000004_4144),
    .const_fix_32_0_1__0000000000000004_4172 (_dup827_const_fix_32_0_1__0000000000000004_4172),
    .const_fix_32_0_1__0000000000000004_4208 (_dup827_const_fix_32_0_1__0000000000000004_4208),
    .const_fix_32_0_1__0000000000000004_4508 (_dup827_const_fix_32_0_1__0000000000000004_4508),
    .const_fix_32_0_1__0000000000000004_4536 (_dup827_const_fix_32_0_1__0000000000000004_4536),
    .const_fix_32_0_1__0000000000000004_4572 (_dup827_const_fix_32_0_1__0000000000000004_4572)
  );
  ADD_2x1 ADD828 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:974:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL826__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:972:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_706_2583_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2601:146
    ._dfc_wire_100                          (_ADD828__dfc_wire_100)
  );
  MUL_2x1 MUL829 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:975:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_689_2580_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2598:146
    ._dfc_wire_104                          (_dup823__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:969:111
    ._dfc_wire_107                          (_MUL829__dfc_wire_107)
  );
  dup_1x2 dup830 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:976:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD828__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:974:130
    ._dfc_wire_68_105 (_dup830__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup830__dfc_wire_68_113)
  );
  ADD_2x1 ADD831 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:977:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup830__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:976:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_60_2579_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2597:142
    ._dfc_wire_100                          (_ADD831__dfc_wire_100)
  );
  SHR3_1x1 SHR3832 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:978:89
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_ADD831__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:977:130
    ._dfc_wire_1968 (_SHR3832__dfc_wire_1968)
  );
  MUL_2x1 MUL833 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:979:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_692_2577_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2595:146
    ._dfc_wire_104                          (_dup824__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:970:111
    ._dfc_wire_107                          (_MUL833__dfc_wire_107)
  );
  SUB_2x1 SUB834 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:980:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup830__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:976:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_125_2576_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2594:146
    ._dfc_wire_121    (_SUB834__dfc_wire_121)
  );
  SHR3_1x1 SHR3835 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:981:89
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB834__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:980:109
    ._dfc_wire_1968 (_SHR3835__dfc_wire_1968)
  );
  dup_1x2 dup836 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:982:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST817__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:963:84
    ._dfc_wire_68_105 (_dup836__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup836__dfc_wire_68_113)
  );
  dup_1x2 dup837 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:983:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST818__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:964:84
    ._dfc_wire_68_105 (_dup837__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup837__dfc_wire_68_113)
  );
  ADD_2x1 ADD838 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:984:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_28_2570_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2588:142
    .const_fix_32_0_1__0000000000000080_102 (_dup837__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:983:111
    ._dfc_wire_100                          (_ADD838__dfc_wire_100)
  );
  MUL_2x1 MUL839 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:985:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_913_2567_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2585:146
    ._dfc_wire_104                          (_ADD838__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:984:130
    ._dfc_wire_107                          (_MUL839__dfc_wire_107)
  );
  ADD_2x1 ADD840 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:986:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL839__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:985:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_842_2565_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2583:146
    ._dfc_wire_100                          (_ADD840__dfc_wire_100)
  );
  MUL_2x1 MUL841 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:987:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_749_3067_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3085:146
    ._dfc_wire_104                          (_dup836__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:982:111
    ._dfc_wire_107                          (_MUL841__dfc_wire_107)
  );
  dup_1x2 dup842 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:988:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD840__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:986:130
    ._dfc_wire_68_105 (_dup842__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup842__dfc_wire_68_113)
  );
  SUB_2x1 SUB843 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:989:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup842__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:988:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_209_3063_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3081:146
    ._dfc_wire_121    (_SUB843__dfc_wire_121)
  );
  SHR3_1x1 SHR3844 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:990:89
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB843__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:989:109
    ._dfc_wire_1968 (_SHR3844__dfc_wire_1968)
  );
  MUL_2x1 MUL845 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:991:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_835_3057_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3075:146
    ._dfc_wire_104                          (_dup837__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:983:111
    ._dfc_wire_107                          (_MUL845__dfc_wire_107)
  );
  SUB_2x1 SUB846 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:992:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup842__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:988:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_218_3055_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3073:146
    ._dfc_wire_121    (_SUB846__dfc_wire_121)
  );
  SHR3_1x1 SHR3847 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:993:89
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB846__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:992:109
    ._dfc_wire_1968 (_SHR3847__dfc_wire_1968)
  );
  dup_1x2 dup848 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:994:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD822__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:968:130
    ._dfc_wire_68_105 (_dup848__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup848__dfc_wire_68_113)
  );
  dup_1x2 dup849 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:995:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHL8812__dfc_wire_1923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:958:89
    ._dfc_wire_68_105 (_dup849__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup849__dfc_wire_68_113)
  );
  ADD_2x1 ADD850 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:996:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup848__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:994:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_126_3046_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3064:146
    ._dfc_wire_100                          (_ADD850__dfc_wire_100)
  );
  SUB_2x1 SUB851 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:997:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup848__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:994:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_126_3044_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3062:146
    ._dfc_wire_121    (_SUB851__dfc_wire_121)
  );
  dup_1x2 dup852 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:998:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST814__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:960:84
    ._dfc_wire_68_105 (_dup852__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup852__dfc_wire_68_113)
  );
  dup_1x2 dup853 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:999:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST813__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:959:84
    ._dfc_wire_68_105 (_dup853__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup853__dfc_wire_68_113)
  );
  ADD_2x1 ADD854 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1000:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_86_3034_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3052:142
    .const_fix_32_0_1__0000000000000080_102 (_dup853__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:999:111
    ._dfc_wire_100                          (_ADD854__dfc_wire_100)
  );
  MUL_2x1 MUL855 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1001:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_822_3030_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3048:146
    ._dfc_wire_104                          (_ADD854__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1000:130
    ._dfc_wire_107                          (_MUL855__dfc_wire_107)
  );
  ADD_2x1 ADD856 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1002:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL855__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1001:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_741_3230_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3248:146
    ._dfc_wire_100                          (_ADD856__dfc_wire_100)
  );
  MUL_2x1 MUL857 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1003:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_787_3028_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3046:146
    ._dfc_wire_104                          (_dup853__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:999:111
    ._dfc_wire_107                          (_MUL857__dfc_wire_107)
  );
  dup_1x2 dup858 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1004:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD856__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1002:130
    ._dfc_wire_68_105 (_dup858__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup858__dfc_wire_68_113)
  );
  SUB_2x1 SUB859 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1005:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup858__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1004:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_136_3026_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3044:146
    ._dfc_wire_121    (_SUB859__dfc_wire_121)
  );
  SHR3_1x1 SHR3860 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1006:89
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB859__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1005:109
    ._dfc_wire_1968 (_SHR3860__dfc_wire_1968)
  );
  MUL_2x1 MUL861 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1007:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_757_3021_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3039:146
    ._dfc_wire_104                          (_dup852__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:998:111
    ._dfc_wire_107                          (_MUL861__dfc_wire_107)
  );
  ADD_2x1 ADD862 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1008:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup858__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1004:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_159_3018_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3036:146
    ._dfc_wire_100                          (_ADD862__dfc_wire_100)
  );
  SHR3_1x1 SHR3863 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1009:89
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_ADD862__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1008:130
    ._dfc_wire_1968 (_SHR3863__dfc_wire_1968)
  );
  dup_1x2 dup864 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1010:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR3832__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:978:89
    ._dfc_wire_68_105 (_dup864__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup864__dfc_wire_68_113)
  );
  dup_1x2 dup865 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1011:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR3844__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:990:89
    ._dfc_wire_68_105 (_dup865__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup865__dfc_wire_68_113)
  );
  ADD_2x1 ADD866 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1012:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_225_3012_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3030:146
    .const_fix_32_0_1__0000000000000080_102 (_dup865__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1011:111
    ._dfc_wire_100                          (_ADD866__dfc_wire_100)
  );
  SUB_2x1 SUB867 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1013:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_225_3010_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3028:146
    ._dfc_wire_118    (_dup865__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1011:111
    ._dfc_wire_121    (_SUB867__dfc_wire_121)
  );
  dup_1x2 dup868 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1014:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR3835__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:981:89
    ._dfc_wire_68_105 (_dup868__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup868__dfc_wire_68_113)
  );
  dup_1x2 dup869 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1015:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR3847__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:993:89
    ._dfc_wire_68_105 (_dup869__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup869__dfc_wire_68_113)
  );
  ADD_2x1 ADD870 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1016:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_206_3002_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3020:146
    .const_fix_32_0_1__0000000000000080_102 (_dup869__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1015:111
    ._dfc_wire_100                          (_ADD870__dfc_wire_100)
  );
  SUB_2x1 SUB871 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1017:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_206_2998_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3016:146
    ._dfc_wire_118    (_dup869__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1015:111
    ._dfc_wire_121    (_SUB871__dfc_wire_121)
  );
  dup_1x2 dup872 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1018:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD850__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:996:130
    ._dfc_wire_68_105 (_dup872__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup872__dfc_wire_68_113)
  );
  dup_1x2 dup873 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1019:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR3863__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1009:89
    ._dfc_wire_68_105 (_dup873__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup873__dfc_wire_68_113)
  );
  ADD_2x1 ADD874 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1020:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_130_2995_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3013:146
    .const_fix_32_0_1__0000000000000080_102 (_dup873__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1019:111
    ._dfc_wire_100                          (_ADD874__dfc_wire_100)
  );
  SUB_2x1 SUB875 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1021:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_130_3211_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3229:146
    ._dfc_wire_118    (_dup873__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1019:111
    ._dfc_wire_121    (_SUB875__dfc_wire_121)
  );
  dup_1x2 dup876 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1022:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB851__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:997:109
    ._dfc_wire_68_105 (_dup876__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup876__dfc_wire_68_113)
  );
  dup_1x2 dup877 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1023:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR3860__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1006:89
    ._dfc_wire_68_105 (_dup877__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup877__dfc_wire_68_113)
  );
  ADD_2x1 ADD878 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1024:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_99_2992_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3010:142
    .const_fix_32_0_1__0000000000000080_102 (_dup877__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1023:111
    ._dfc_wire_100                          (_ADD878__dfc_wire_100)
  );
  SUB_2x1 SUB879 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1025:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_99_2991_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3009:142
    ._dfc_wire_118    (_dup877__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1023:111
    ._dfc_wire_121    (_SUB879__dfc_wire_121)
  );
  dup_1x2 dup880 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1026:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB867__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1013:109
    ._dfc_wire_68_105 (_dup880__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup880__dfc_wire_68_113)
  );
  dup_1x2 dup881 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1027:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB871__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1017:109
    ._dfc_wire_68_105 (_dup881__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup881__dfc_wire_68_113)
  );
  ADD_2x1 ADD882 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1028:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup880__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1026:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_6_2987_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3005:138
    ._dfc_wire_100                          (_ADD882__dfc_wire_100)
  );
  MUL_2x1 MUL883 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1029:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1404_2986_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3004:150
    ._dfc_wire_104                          (_ADD882__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1028:130
    ._dfc_wire_107                          (_MUL883__dfc_wire_107)
  );
  ADD_2x1 ADD884 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1030:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL883__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1029:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1557_2983_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3001:150
    ._dfc_wire_100                          (_ADD884__dfc_wire_100)
  );
  SHR8_1x1 SHR8885 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1031:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD884__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1030:130
    ._dfc_wire_216 (_SHR8885__dfc_wire_216)
  );
  SUB_2x1 SUB886 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1032:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup880__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1026:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_6_2981_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2999:138
    ._dfc_wire_121    (_SUB886__dfc_wire_121)
  );
  MUL_2x1 MUL887 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1033:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1391_2980_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2998:150
    ._dfc_wire_104                          (_SUB886__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1032:109
    ._dfc_wire_107                          (_MUL887__dfc_wire_107)
  );
  ADD_2x1 ADD888 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1034:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL887__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1033:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1564_2979_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2997:150
    ._dfc_wire_100                          (_ADD888__dfc_wire_100)
  );
  SHR8_1x1 SHR8889 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1035:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD888__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1034:130
    ._dfc_wire_216 (_SHR8889__dfc_wire_216)
  );
  dup_1x2 dup890 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1036:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD874__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1020:130
    ._dfc_wire_68_105 (_dup890__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup890__dfc_wire_68_113)
  );
  dup_1x2 dup891 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1037:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD866__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1012:130
    ._dfc_wire_68_105 (_dup891__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup891__dfc_wire_68_113)
  );
  ADD_2x1 ADD892 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1038:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_190_2978_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2996:146
    .const_fix_32_0_1__0000000000000080_102 (_dup891__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1037:111
    ._dfc_wire_100                          (_ADD892__dfc_wire_100)
  );
  SHR14_1x1 SHR14893 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1039:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD892__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1038:130
    ._dfc_wire_2103 (_SHR14893__dfc_wire_2103)
  );
  dup_1x3 dup894 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1040:148
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR14893__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1039:93
    ._dfc_wire_2103_2106 (_dup894__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup894__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup894__dfc_wire_2103_2113)
  );
  dup_1x128 dup895 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .clock                                   (clock),
    .reset                                   (reset),
    .const_fix_32_0_1__00000000000000ff      (_const2146_const_fix_32_0_1__00000000000000ff),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2166:90
    .const_fix_32_0_1__00000000000000ff_2107 (_dup895_const_fix_32_0_1__00000000000000ff_2107),
    .const_fix_32_0_1__00000000000000ff_2111 (_dup895_const_fix_32_0_1__00000000000000ff_2111),
    .const_fix_32_0_1__00000000000000ff_2129 (_dup895_const_fix_32_0_1__00000000000000ff_2129),
    .const_fix_32_0_1__00000000000000ff_2133 (_dup895_const_fix_32_0_1__00000000000000ff_2133),
    .const_fix_32_0_1__00000000000000ff_2151 (_dup895_const_fix_32_0_1__00000000000000ff_2151),
    .const_fix_32_0_1__00000000000000ff_2155 (_dup895_const_fix_32_0_1__00000000000000ff_2155),
    .const_fix_32_0_1__00000000000000ff_2173 (_dup895_const_fix_32_0_1__00000000000000ff_2173),
    .const_fix_32_0_1__00000000000000ff_2177 (_dup895_const_fix_32_0_1__00000000000000ff_2177),
    .const_fix_32_0_1__00000000000000ff_2195 (_dup895_const_fix_32_0_1__00000000000000ff_2195),
    .const_fix_32_0_1__00000000000000ff_2199 (_dup895_const_fix_32_0_1__00000000000000ff_2199),
    .const_fix_32_0_1__00000000000000ff_2217 (_dup895_const_fix_32_0_1__00000000000000ff_2217),
    .const_fix_32_0_1__00000000000000ff_2221 (_dup895_const_fix_32_0_1__00000000000000ff_2221),
    .const_fix_32_0_1__00000000000000ff_2239 (_dup895_const_fix_32_0_1__00000000000000ff_2239),
    .const_fix_32_0_1__00000000000000ff_2243 (_dup895_const_fix_32_0_1__00000000000000ff_2243),
    .const_fix_32_0_1__00000000000000ff_2261 (_dup895_const_fix_32_0_1__00000000000000ff_2261),
    .const_fix_32_0_1__00000000000000ff_2265 (_dup895_const_fix_32_0_1__00000000000000ff_2265),
    .const_fix_32_0_1__00000000000000ff_2471 (_dup895_const_fix_32_0_1__00000000000000ff_2471),
    .const_fix_32_0_1__00000000000000ff_2475 (_dup895_const_fix_32_0_1__00000000000000ff_2475),
    .const_fix_32_0_1__00000000000000ff_2493 (_dup895_const_fix_32_0_1__00000000000000ff_2493),
    .const_fix_32_0_1__00000000000000ff_2497 (_dup895_const_fix_32_0_1__00000000000000ff_2497),
    .const_fix_32_0_1__00000000000000ff_2515 (_dup895_const_fix_32_0_1__00000000000000ff_2515),
    .const_fix_32_0_1__00000000000000ff_2519 (_dup895_const_fix_32_0_1__00000000000000ff_2519),
    .const_fix_32_0_1__00000000000000ff_2537 (_dup895_const_fix_32_0_1__00000000000000ff_2537),
    .const_fix_32_0_1__00000000000000ff_2541 (_dup895_const_fix_32_0_1__00000000000000ff_2541),
    .const_fix_32_0_1__00000000000000ff_2559 (_dup895_const_fix_32_0_1__00000000000000ff_2559),
    .const_fix_32_0_1__00000000000000ff_2563 (_dup895_const_fix_32_0_1__00000000000000ff_2563),
    .const_fix_32_0_1__00000000000000ff_2581 (_dup895_const_fix_32_0_1__00000000000000ff_2581),
    .const_fix_32_0_1__00000000000000ff_2585 (_dup895_const_fix_32_0_1__00000000000000ff_2585),
    .const_fix_32_0_1__00000000000000ff_2603 (_dup895_const_fix_32_0_1__00000000000000ff_2603),
    .const_fix_32_0_1__00000000000000ff_2607 (_dup895_const_fix_32_0_1__00000000000000ff_2607),
    .const_fix_32_0_1__00000000000000ff_2625 (_dup895_const_fix_32_0_1__00000000000000ff_2625),
    .const_fix_32_0_1__00000000000000ff_2629 (_dup895_const_fix_32_0_1__00000000000000ff_2629),
    .const_fix_32_0_1__00000000000000ff_2835 (_dup895_const_fix_32_0_1__00000000000000ff_2835),
    .const_fix_32_0_1__00000000000000ff_2839 (_dup895_const_fix_32_0_1__00000000000000ff_2839),
    .const_fix_32_0_1__00000000000000ff_2857 (_dup895_const_fix_32_0_1__00000000000000ff_2857),
    .const_fix_32_0_1__00000000000000ff_2861 (_dup895_const_fix_32_0_1__00000000000000ff_2861),
    .const_fix_32_0_1__00000000000000ff_2879 (_dup895_const_fix_32_0_1__00000000000000ff_2879),
    .const_fix_32_0_1__00000000000000ff_2883 (_dup895_const_fix_32_0_1__00000000000000ff_2883),
    .const_fix_32_0_1__00000000000000ff_2901 (_dup895_const_fix_32_0_1__00000000000000ff_2901),
    .const_fix_32_0_1__00000000000000ff_2905 (_dup895_const_fix_32_0_1__00000000000000ff_2905),
    .const_fix_32_0_1__00000000000000ff_2923 (_dup895_const_fix_32_0_1__00000000000000ff_2923),
    .const_fix_32_0_1__00000000000000ff_2927 (_dup895_const_fix_32_0_1__00000000000000ff_2927),
    .const_fix_32_0_1__00000000000000ff_2945 (_dup895_const_fix_32_0_1__00000000000000ff_2945),
    .const_fix_32_0_1__00000000000000ff_2949 (_dup895_const_fix_32_0_1__00000000000000ff_2949),
    .const_fix_32_0_1__00000000000000ff_2967 (_dup895_const_fix_32_0_1__00000000000000ff_2967),
    .const_fix_32_0_1__00000000000000ff_2971 (_dup895_const_fix_32_0_1__00000000000000ff_2971),
    .const_fix_32_0_1__00000000000000ff_2989 (_dup895_const_fix_32_0_1__00000000000000ff_2989),
    .const_fix_32_0_1__00000000000000ff_2993 (_dup895_const_fix_32_0_1__00000000000000ff_2993),
    .const_fix_32_0_1__00000000000000ff_3199 (_dup895_const_fix_32_0_1__00000000000000ff_3199),
    .const_fix_32_0_1__00000000000000ff_3203 (_dup895_const_fix_32_0_1__00000000000000ff_3203),
    .const_fix_32_0_1__00000000000000ff_3221 (_dup895_const_fix_32_0_1__00000000000000ff_3221),
    .const_fix_32_0_1__00000000000000ff_3225 (_dup895_const_fix_32_0_1__00000000000000ff_3225),
    .const_fix_32_0_1__00000000000000ff_3243 (_dup895_const_fix_32_0_1__00000000000000ff_3243),
    .const_fix_32_0_1__00000000000000ff_3247 (_dup895_const_fix_32_0_1__00000000000000ff_3247),
    .const_fix_32_0_1__00000000000000ff_3265 (_dup895_const_fix_32_0_1__00000000000000ff_3265),
    .const_fix_32_0_1__00000000000000ff_3269 (_dup895_const_fix_32_0_1__00000000000000ff_3269),
    .const_fix_32_0_1__00000000000000ff_3287 (_dup895_const_fix_32_0_1__00000000000000ff_3287),
    .const_fix_32_0_1__00000000000000ff_3291 (_dup895_const_fix_32_0_1__00000000000000ff_3291),
    .const_fix_32_0_1__00000000000000ff_3309 (_dup895_const_fix_32_0_1__00000000000000ff_3309),
    .const_fix_32_0_1__00000000000000ff_3313 (_dup895_const_fix_32_0_1__00000000000000ff_3313),
    .const_fix_32_0_1__00000000000000ff_3331 (_dup895_const_fix_32_0_1__00000000000000ff_3331),
    .const_fix_32_0_1__00000000000000ff_3335 (_dup895_const_fix_32_0_1__00000000000000ff_3335),
    .const_fix_32_0_1__00000000000000ff_3353 (_dup895_const_fix_32_0_1__00000000000000ff_3353),
    .const_fix_32_0_1__00000000000000ff_3357 (_dup895_const_fix_32_0_1__00000000000000ff_3357),
    .const_fix_32_0_1__00000000000000ff_3563 (_dup895_const_fix_32_0_1__00000000000000ff_3563),
    .const_fix_32_0_1__00000000000000ff_3567 (_dup895_const_fix_32_0_1__00000000000000ff_3567),
    .const_fix_32_0_1__00000000000000ff_3585 (_dup895_const_fix_32_0_1__00000000000000ff_3585),
    .const_fix_32_0_1__00000000000000ff_3589 (_dup895_const_fix_32_0_1__00000000000000ff_3589),
    .const_fix_32_0_1__00000000000000ff_3607 (_dup895_const_fix_32_0_1__00000000000000ff_3607),
    .const_fix_32_0_1__00000000000000ff_3611 (_dup895_const_fix_32_0_1__00000000000000ff_3611),
    .const_fix_32_0_1__00000000000000ff_3629 (_dup895_const_fix_32_0_1__00000000000000ff_3629),
    .const_fix_32_0_1__00000000000000ff_3633 (_dup895_const_fix_32_0_1__00000000000000ff_3633),
    .const_fix_32_0_1__00000000000000ff_3651 (_dup895_const_fix_32_0_1__00000000000000ff_3651),
    .const_fix_32_0_1__00000000000000ff_3655 (_dup895_const_fix_32_0_1__00000000000000ff_3655),
    .const_fix_32_0_1__00000000000000ff_3673 (_dup895_const_fix_32_0_1__00000000000000ff_3673),
    .const_fix_32_0_1__00000000000000ff_3677 (_dup895_const_fix_32_0_1__00000000000000ff_3677),
    .const_fix_32_0_1__00000000000000ff_3695 (_dup895_const_fix_32_0_1__00000000000000ff_3695),
    .const_fix_32_0_1__00000000000000ff_3699 (_dup895_const_fix_32_0_1__00000000000000ff_3699),
    .const_fix_32_0_1__00000000000000ff_3717 (_dup895_const_fix_32_0_1__00000000000000ff_3717),
    .const_fix_32_0_1__00000000000000ff_3721 (_dup895_const_fix_32_0_1__00000000000000ff_3721),
    .const_fix_32_0_1__00000000000000ff_3927 (_dup895_const_fix_32_0_1__00000000000000ff_3927),
    .const_fix_32_0_1__00000000000000ff_3931 (_dup895_const_fix_32_0_1__00000000000000ff_3931),
    .const_fix_32_0_1__00000000000000ff_3949 (_dup895_const_fix_32_0_1__00000000000000ff_3949),
    .const_fix_32_0_1__00000000000000ff_3953 (_dup895_const_fix_32_0_1__00000000000000ff_3953),
    .const_fix_32_0_1__00000000000000ff_3971 (_dup895_const_fix_32_0_1__00000000000000ff_3971),
    .const_fix_32_0_1__00000000000000ff_3975 (_dup895_const_fix_32_0_1__00000000000000ff_3975),
    .const_fix_32_0_1__00000000000000ff_3993 (_dup895_const_fix_32_0_1__00000000000000ff_3993),
    .const_fix_32_0_1__00000000000000ff_3997 (_dup895_const_fix_32_0_1__00000000000000ff_3997),
    .const_fix_32_0_1__00000000000000ff_4015 (_dup895_const_fix_32_0_1__00000000000000ff_4015),
    .const_fix_32_0_1__00000000000000ff_4019 (_dup895_const_fix_32_0_1__00000000000000ff_4019),
    .const_fix_32_0_1__00000000000000ff_4037 (_dup895_const_fix_32_0_1__00000000000000ff_4037),
    .const_fix_32_0_1__00000000000000ff_4041 (_dup895_const_fix_32_0_1__00000000000000ff_4041),
    .const_fix_32_0_1__00000000000000ff_4059 (_dup895_const_fix_32_0_1__00000000000000ff_4059),
    .const_fix_32_0_1__00000000000000ff_4063 (_dup895_const_fix_32_0_1__00000000000000ff_4063),
    .const_fix_32_0_1__00000000000000ff_4081 (_dup895_const_fix_32_0_1__00000000000000ff_4081),
    .const_fix_32_0_1__00000000000000ff_4085 (_dup895_const_fix_32_0_1__00000000000000ff_4085),
    .const_fix_32_0_1__00000000000000ff_4291 (_dup895_const_fix_32_0_1__00000000000000ff_4291),
    .const_fix_32_0_1__00000000000000ff_4295 (_dup895_const_fix_32_0_1__00000000000000ff_4295),
    .const_fix_32_0_1__00000000000000ff_4313 (_dup895_const_fix_32_0_1__00000000000000ff_4313),
    .const_fix_32_0_1__00000000000000ff_4317 (_dup895_const_fix_32_0_1__00000000000000ff_4317),
    .const_fix_32_0_1__00000000000000ff_4335 (_dup895_const_fix_32_0_1__00000000000000ff_4335),
    .const_fix_32_0_1__00000000000000ff_4339 (_dup895_const_fix_32_0_1__00000000000000ff_4339),
    .const_fix_32_0_1__00000000000000ff_4357 (_dup895_const_fix_32_0_1__00000000000000ff_4357),
    .const_fix_32_0_1__00000000000000ff_4361 (_dup895_const_fix_32_0_1__00000000000000ff_4361),
    .const_fix_32_0_1__00000000000000ff_4379 (_dup895_const_fix_32_0_1__00000000000000ff_4379),
    .const_fix_32_0_1__00000000000000ff_4383 (_dup895_const_fix_32_0_1__00000000000000ff_4383),
    .const_fix_32_0_1__00000000000000ff_4401 (_dup895_const_fix_32_0_1__00000000000000ff_4401),
    .const_fix_32_0_1__00000000000000ff_4405 (_dup895_const_fix_32_0_1__00000000000000ff_4405),
    .const_fix_32_0_1__00000000000000ff_4423 (_dup895_const_fix_32_0_1__00000000000000ff_4423),
    .const_fix_32_0_1__00000000000000ff_4427 (_dup895_const_fix_32_0_1__00000000000000ff_4427),
    .const_fix_32_0_1__00000000000000ff_4445 (_dup895_const_fix_32_0_1__00000000000000ff_4445),
    .const_fix_32_0_1__00000000000000ff_4449 (_dup895_const_fix_32_0_1__00000000000000ff_4449),
    .const_fix_32_0_1__00000000000000ff_4655 (_dup895_const_fix_32_0_1__00000000000000ff_4655),
    .const_fix_32_0_1__00000000000000ff_4659 (_dup895_const_fix_32_0_1__00000000000000ff_4659),
    .const_fix_32_0_1__00000000000000ff_4677 (_dup895_const_fix_32_0_1__00000000000000ff_4677),
    .const_fix_32_0_1__00000000000000ff_4681 (_dup895_const_fix_32_0_1__00000000000000ff_4681),
    .const_fix_32_0_1__00000000000000ff_4699 (_dup895_const_fix_32_0_1__00000000000000ff_4699),
    .const_fix_32_0_1__00000000000000ff_4703 (_dup895_const_fix_32_0_1__00000000000000ff_4703),
    .const_fix_32_0_1__00000000000000ff_4721 (_dup895_const_fix_32_0_1__00000000000000ff_4721),
    .const_fix_32_0_1__00000000000000ff_4725 (_dup895_const_fix_32_0_1__00000000000000ff_4725),
    .const_fix_32_0_1__00000000000000ff_4743 (_dup895_const_fix_32_0_1__00000000000000ff_4743),
    .const_fix_32_0_1__00000000000000ff_4747 (_dup895_const_fix_32_0_1__00000000000000ff_4747),
    .const_fix_32_0_1__00000000000000ff_4765 (_dup895_const_fix_32_0_1__00000000000000ff_4765),
    .const_fix_32_0_1__00000000000000ff_4769 (_dup895_const_fix_32_0_1__00000000000000ff_4769),
    .const_fix_32_0_1__00000000000000ff_4787 (_dup895_const_fix_32_0_1__00000000000000ff_4787),
    .const_fix_32_0_1__00000000000000ff_4791 (_dup895_const_fix_32_0_1__00000000000000ff_4791),
    .const_fix_32_0_1__00000000000000ff_4809 (_dup895_const_fix_32_0_1__00000000000000ff_4809),
    .const_fix_32_0_1__00000000000000ff_4813 (_dup895_const_fix_32_0_1__00000000000000ff_4813)
  );
  GT_2x1 GT896 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1042:134
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup894__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1040:148
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1560_2721_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2739:150
    ._dfc_wire_2105                          (_GT896__dfc_wire_2105)
  );
  MUX_3x1 MUX897 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1043:163
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT896__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1042:134
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_40_2718_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2736:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1600_2719_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2737:150
    ._dfc_wire_2108                          (_MUX897__dfc_wire_2108)
  );
  dup_1x128 dup898 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .clock                                   (clock),
    .reset                                   (reset),
    .const_fix_32_0_1__00000000000000ff      (_const2086_const_fix_32_0_1__ffffffffffffff00),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2159:90
    .const_fix_32_0_1__00000000000000ff_2107 (_dup898_const_fix_32_0_1__00000000000000ff_2107),
    .const_fix_32_0_1__00000000000000ff_2111 (_dup898_const_fix_32_0_1__00000000000000ff_2111),
    .const_fix_32_0_1__00000000000000ff_2129 (_dup898_const_fix_32_0_1__00000000000000ff_2129),
    .const_fix_32_0_1__00000000000000ff_2133 (_dup898_const_fix_32_0_1__00000000000000ff_2133),
    .const_fix_32_0_1__00000000000000ff_2151 (_dup898_const_fix_32_0_1__00000000000000ff_2151),
    .const_fix_32_0_1__00000000000000ff_2155 (_dup898_const_fix_32_0_1__00000000000000ff_2155),
    .const_fix_32_0_1__00000000000000ff_2173 (_dup898_const_fix_32_0_1__00000000000000ff_2173),
    .const_fix_32_0_1__00000000000000ff_2177 (_dup898_const_fix_32_0_1__00000000000000ff_2177),
    .const_fix_32_0_1__00000000000000ff_2195 (_dup898_const_fix_32_0_1__00000000000000ff_2195),
    .const_fix_32_0_1__00000000000000ff_2199 (_dup898_const_fix_32_0_1__00000000000000ff_2199),
    .const_fix_32_0_1__00000000000000ff_2217 (_dup898_const_fix_32_0_1__00000000000000ff_2217),
    .const_fix_32_0_1__00000000000000ff_2221 (_dup898_const_fix_32_0_1__00000000000000ff_2221),
    .const_fix_32_0_1__00000000000000ff_2239 (_dup898_const_fix_32_0_1__00000000000000ff_2239),
    .const_fix_32_0_1__00000000000000ff_2243 (_dup898_const_fix_32_0_1__00000000000000ff_2243),
    .const_fix_32_0_1__00000000000000ff_2261 (_dup898_const_fix_32_0_1__00000000000000ff_2261),
    .const_fix_32_0_1__00000000000000ff_2265 (_dup898_const_fix_32_0_1__00000000000000ff_2265),
    .const_fix_32_0_1__00000000000000ff_2471 (_dup898_const_fix_32_0_1__00000000000000ff_2471),
    .const_fix_32_0_1__00000000000000ff_2475 (_dup898_const_fix_32_0_1__00000000000000ff_2475),
    .const_fix_32_0_1__00000000000000ff_2493 (_dup898_const_fix_32_0_1__00000000000000ff_2493),
    .const_fix_32_0_1__00000000000000ff_2497 (_dup898_const_fix_32_0_1__00000000000000ff_2497),
    .const_fix_32_0_1__00000000000000ff_2515 (_dup898_const_fix_32_0_1__00000000000000ff_2515),
    .const_fix_32_0_1__00000000000000ff_2519 (_dup898_const_fix_32_0_1__00000000000000ff_2519),
    .const_fix_32_0_1__00000000000000ff_2537 (_dup898_const_fix_32_0_1__00000000000000ff_2537),
    .const_fix_32_0_1__00000000000000ff_2541 (_dup898_const_fix_32_0_1__00000000000000ff_2541),
    .const_fix_32_0_1__00000000000000ff_2559 (_dup898_const_fix_32_0_1__00000000000000ff_2559),
    .const_fix_32_0_1__00000000000000ff_2563 (_dup898_const_fix_32_0_1__00000000000000ff_2563),
    .const_fix_32_0_1__00000000000000ff_2581 (_dup898_const_fix_32_0_1__00000000000000ff_2581),
    .const_fix_32_0_1__00000000000000ff_2585 (_dup898_const_fix_32_0_1__00000000000000ff_2585),
    .const_fix_32_0_1__00000000000000ff_2603 (_dup898_const_fix_32_0_1__00000000000000ff_2603),
    .const_fix_32_0_1__00000000000000ff_2607 (_dup898_const_fix_32_0_1__00000000000000ff_2607),
    .const_fix_32_0_1__00000000000000ff_2625 (_dup898_const_fix_32_0_1__00000000000000ff_2625),
    .const_fix_32_0_1__00000000000000ff_2629 (_dup898_const_fix_32_0_1__00000000000000ff_2629),
    .const_fix_32_0_1__00000000000000ff_2835 (_dup898_const_fix_32_0_1__00000000000000ff_2835),
    .const_fix_32_0_1__00000000000000ff_2839 (_dup898_const_fix_32_0_1__00000000000000ff_2839),
    .const_fix_32_0_1__00000000000000ff_2857 (_dup898_const_fix_32_0_1__00000000000000ff_2857),
    .const_fix_32_0_1__00000000000000ff_2861 (_dup898_const_fix_32_0_1__00000000000000ff_2861),
    .const_fix_32_0_1__00000000000000ff_2879 (_dup898_const_fix_32_0_1__00000000000000ff_2879),
    .const_fix_32_0_1__00000000000000ff_2883 (_dup898_const_fix_32_0_1__00000000000000ff_2883),
    .const_fix_32_0_1__00000000000000ff_2901 (_dup898_const_fix_32_0_1__00000000000000ff_2901),
    .const_fix_32_0_1__00000000000000ff_2905 (_dup898_const_fix_32_0_1__00000000000000ff_2905),
    .const_fix_32_0_1__00000000000000ff_2923 (_dup898_const_fix_32_0_1__00000000000000ff_2923),
    .const_fix_32_0_1__00000000000000ff_2927 (_dup898_const_fix_32_0_1__00000000000000ff_2927),
    .const_fix_32_0_1__00000000000000ff_2945 (_dup898_const_fix_32_0_1__00000000000000ff_2945),
    .const_fix_32_0_1__00000000000000ff_2949 (_dup898_const_fix_32_0_1__00000000000000ff_2949),
    .const_fix_32_0_1__00000000000000ff_2967 (_dup898_const_fix_32_0_1__00000000000000ff_2967),
    .const_fix_32_0_1__00000000000000ff_2971 (_dup898_const_fix_32_0_1__00000000000000ff_2971),
    .const_fix_32_0_1__00000000000000ff_2989 (_dup898_const_fix_32_0_1__00000000000000ff_2989),
    .const_fix_32_0_1__00000000000000ff_2993 (_dup898_const_fix_32_0_1__00000000000000ff_2993),
    .const_fix_32_0_1__00000000000000ff_3199 (_dup898_const_fix_32_0_1__00000000000000ff_3199),
    .const_fix_32_0_1__00000000000000ff_3203 (_dup898_const_fix_32_0_1__00000000000000ff_3203),
    .const_fix_32_0_1__00000000000000ff_3221 (_dup898_const_fix_32_0_1__00000000000000ff_3221),
    .const_fix_32_0_1__00000000000000ff_3225 (_dup898_const_fix_32_0_1__00000000000000ff_3225),
    .const_fix_32_0_1__00000000000000ff_3243 (_dup898_const_fix_32_0_1__00000000000000ff_3243),
    .const_fix_32_0_1__00000000000000ff_3247 (_dup898_const_fix_32_0_1__00000000000000ff_3247),
    .const_fix_32_0_1__00000000000000ff_3265 (_dup898_const_fix_32_0_1__00000000000000ff_3265),
    .const_fix_32_0_1__00000000000000ff_3269 (_dup898_const_fix_32_0_1__00000000000000ff_3269),
    .const_fix_32_0_1__00000000000000ff_3287 (_dup898_const_fix_32_0_1__00000000000000ff_3287),
    .const_fix_32_0_1__00000000000000ff_3291 (_dup898_const_fix_32_0_1__00000000000000ff_3291),
    .const_fix_32_0_1__00000000000000ff_3309 (_dup898_const_fix_32_0_1__00000000000000ff_3309),
    .const_fix_32_0_1__00000000000000ff_3313 (_dup898_const_fix_32_0_1__00000000000000ff_3313),
    .const_fix_32_0_1__00000000000000ff_3331 (_dup898_const_fix_32_0_1__00000000000000ff_3331),
    .const_fix_32_0_1__00000000000000ff_3335 (_dup898_const_fix_32_0_1__00000000000000ff_3335),
    .const_fix_32_0_1__00000000000000ff_3353 (_dup898_const_fix_32_0_1__00000000000000ff_3353),
    .const_fix_32_0_1__00000000000000ff_3357 (_dup898_const_fix_32_0_1__00000000000000ff_3357),
    .const_fix_32_0_1__00000000000000ff_3563 (_dup898_const_fix_32_0_1__00000000000000ff_3563),
    .const_fix_32_0_1__00000000000000ff_3567 (_dup898_const_fix_32_0_1__00000000000000ff_3567),
    .const_fix_32_0_1__00000000000000ff_3585 (_dup898_const_fix_32_0_1__00000000000000ff_3585),
    .const_fix_32_0_1__00000000000000ff_3589 (_dup898_const_fix_32_0_1__00000000000000ff_3589),
    .const_fix_32_0_1__00000000000000ff_3607 (_dup898_const_fix_32_0_1__00000000000000ff_3607),
    .const_fix_32_0_1__00000000000000ff_3611 (_dup898_const_fix_32_0_1__00000000000000ff_3611),
    .const_fix_32_0_1__00000000000000ff_3629 (_dup898_const_fix_32_0_1__00000000000000ff_3629),
    .const_fix_32_0_1__00000000000000ff_3633 (_dup898_const_fix_32_0_1__00000000000000ff_3633),
    .const_fix_32_0_1__00000000000000ff_3651 (_dup898_const_fix_32_0_1__00000000000000ff_3651),
    .const_fix_32_0_1__00000000000000ff_3655 (_dup898_const_fix_32_0_1__00000000000000ff_3655),
    .const_fix_32_0_1__00000000000000ff_3673 (_dup898_const_fix_32_0_1__00000000000000ff_3673),
    .const_fix_32_0_1__00000000000000ff_3677 (_dup898_const_fix_32_0_1__00000000000000ff_3677),
    .const_fix_32_0_1__00000000000000ff_3695 (_dup898_const_fix_32_0_1__00000000000000ff_3695),
    .const_fix_32_0_1__00000000000000ff_3699 (_dup898_const_fix_32_0_1__00000000000000ff_3699),
    .const_fix_32_0_1__00000000000000ff_3717 (_dup898_const_fix_32_0_1__00000000000000ff_3717),
    .const_fix_32_0_1__00000000000000ff_3721 (_dup898_const_fix_32_0_1__00000000000000ff_3721),
    .const_fix_32_0_1__00000000000000ff_3927 (_dup898_const_fix_32_0_1__00000000000000ff_3927),
    .const_fix_32_0_1__00000000000000ff_3931 (_dup898_const_fix_32_0_1__00000000000000ff_3931),
    .const_fix_32_0_1__00000000000000ff_3949 (_dup898_const_fix_32_0_1__00000000000000ff_3949),
    .const_fix_32_0_1__00000000000000ff_3953 (_dup898_const_fix_32_0_1__00000000000000ff_3953),
    .const_fix_32_0_1__00000000000000ff_3971 (_dup898_const_fix_32_0_1__00000000000000ff_3971),
    .const_fix_32_0_1__00000000000000ff_3975 (_dup898_const_fix_32_0_1__00000000000000ff_3975),
    .const_fix_32_0_1__00000000000000ff_3993 (_dup898_const_fix_32_0_1__00000000000000ff_3993),
    .const_fix_32_0_1__00000000000000ff_3997 (_dup898_const_fix_32_0_1__00000000000000ff_3997),
    .const_fix_32_0_1__00000000000000ff_4015 (_dup898_const_fix_32_0_1__00000000000000ff_4015),
    .const_fix_32_0_1__00000000000000ff_4019 (_dup898_const_fix_32_0_1__00000000000000ff_4019),
    .const_fix_32_0_1__00000000000000ff_4037 (_dup898_const_fix_32_0_1__00000000000000ff_4037),
    .const_fix_32_0_1__00000000000000ff_4041 (_dup898_const_fix_32_0_1__00000000000000ff_4041),
    .const_fix_32_0_1__00000000000000ff_4059 (_dup898_const_fix_32_0_1__00000000000000ff_4059),
    .const_fix_32_0_1__00000000000000ff_4063 (_dup898_const_fix_32_0_1__00000000000000ff_4063),
    .const_fix_32_0_1__00000000000000ff_4081 (_dup898_const_fix_32_0_1__00000000000000ff_4081),
    .const_fix_32_0_1__00000000000000ff_4085 (_dup898_const_fix_32_0_1__00000000000000ff_4085),
    .const_fix_32_0_1__00000000000000ff_4291 (_dup898_const_fix_32_0_1__00000000000000ff_4291),
    .const_fix_32_0_1__00000000000000ff_4295 (_dup898_const_fix_32_0_1__00000000000000ff_4295),
    .const_fix_32_0_1__00000000000000ff_4313 (_dup898_const_fix_32_0_1__00000000000000ff_4313),
    .const_fix_32_0_1__00000000000000ff_4317 (_dup898_const_fix_32_0_1__00000000000000ff_4317),
    .const_fix_32_0_1__00000000000000ff_4335 (_dup898_const_fix_32_0_1__00000000000000ff_4335),
    .const_fix_32_0_1__00000000000000ff_4339 (_dup898_const_fix_32_0_1__00000000000000ff_4339),
    .const_fix_32_0_1__00000000000000ff_4357 (_dup898_const_fix_32_0_1__00000000000000ff_4357),
    .const_fix_32_0_1__00000000000000ff_4361 (_dup898_const_fix_32_0_1__00000000000000ff_4361),
    .const_fix_32_0_1__00000000000000ff_4379 (_dup898_const_fix_32_0_1__00000000000000ff_4379),
    .const_fix_32_0_1__00000000000000ff_4383 (_dup898_const_fix_32_0_1__00000000000000ff_4383),
    .const_fix_32_0_1__00000000000000ff_4401 (_dup898_const_fix_32_0_1__00000000000000ff_4401),
    .const_fix_32_0_1__00000000000000ff_4405 (_dup898_const_fix_32_0_1__00000000000000ff_4405),
    .const_fix_32_0_1__00000000000000ff_4423 (_dup898_const_fix_32_0_1__00000000000000ff_4423),
    .const_fix_32_0_1__00000000000000ff_4427 (_dup898_const_fix_32_0_1__00000000000000ff_4427),
    .const_fix_32_0_1__00000000000000ff_4445 (_dup898_const_fix_32_0_1__00000000000000ff_4445),
    .const_fix_32_0_1__00000000000000ff_4449 (_dup898_const_fix_32_0_1__00000000000000ff_4449),
    .const_fix_32_0_1__00000000000000ff_4655 (_dup898_const_fix_32_0_1__00000000000000ff_4655),
    .const_fix_32_0_1__00000000000000ff_4659 (_dup898_const_fix_32_0_1__00000000000000ff_4659),
    .const_fix_32_0_1__00000000000000ff_4677 (_dup898_const_fix_32_0_1__00000000000000ff_4677),
    .const_fix_32_0_1__00000000000000ff_4681 (_dup898_const_fix_32_0_1__00000000000000ff_4681),
    .const_fix_32_0_1__00000000000000ff_4699 (_dup898_const_fix_32_0_1__00000000000000ff_4699),
    .const_fix_32_0_1__00000000000000ff_4703 (_dup898_const_fix_32_0_1__00000000000000ff_4703),
    .const_fix_32_0_1__00000000000000ff_4721 (_dup898_const_fix_32_0_1__00000000000000ff_4721),
    .const_fix_32_0_1__00000000000000ff_4725 (_dup898_const_fix_32_0_1__00000000000000ff_4725),
    .const_fix_32_0_1__00000000000000ff_4743 (_dup898_const_fix_32_0_1__00000000000000ff_4743),
    .const_fix_32_0_1__00000000000000ff_4747 (_dup898_const_fix_32_0_1__00000000000000ff_4747),
    .const_fix_32_0_1__00000000000000ff_4765 (_dup898_const_fix_32_0_1__00000000000000ff_4765),
    .const_fix_32_0_1__00000000000000ff_4769 (_dup898_const_fix_32_0_1__00000000000000ff_4769),
    .const_fix_32_0_1__00000000000000ff_4787 (_dup898_const_fix_32_0_1__00000000000000ff_4787),
    .const_fix_32_0_1__00000000000000ff_4791 (_dup898_const_fix_32_0_1__00000000000000ff_4791),
    .const_fix_32_0_1__00000000000000ff_4809 (_dup898_const_fix_32_0_1__00000000000000ff_4809),
    .const_fix_32_0_1__00000000000000ff_4813 (_dup898_const_fix_32_0_1__00000000000000ff_4813)
  );
  LT_2x1 LT899 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1045:134
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup894__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1040:148
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1526_2715_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2733:150
    ._dfc_wire_2112                          (_LT899__dfc_wire_2112)
  );
  MUX_3x1 MUX900 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1046:163
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_LT899__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1045:134
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_53_2712_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2730:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1623_2713_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2731:150
    ._dfc_wire_2108                          (_MUX900__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST901 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1047:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX900__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1046:163
    ._dfc_wire_236 (sink__dfc_wire_2119__dfc_wire_4799)
  );
  dup_1x2 dup902 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1048:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD878__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1024:130
    ._dfc_wire_68_105 (_dup902__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup902__dfc_wire_68_113)
  );
  dup_1x2 dup903 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1049:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR8885__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1031:87
    ._dfc_wire_68_105 (_dup903__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup903__dfc_wire_68_113)
  );
  ADD_2x1 ADD904 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1050:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_460_2707_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2725:146
    .const_fix_32_0_1__0000000000000080_102 (_dup903__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1049:111
    ._dfc_wire_100                          (_ADD904__dfc_wire_100)
  );
  SHR14_1x1 SHR14905 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1051:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD904__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1050:130
    ._dfc_wire_2103 (_SHR14905__dfc_wire_2103)
  );
  dup_1x3 dup906 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1052:148
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR14905__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1051:93
    ._dfc_wire_2103_2106 (_dup906__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup906__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup906__dfc_wire_2103_2113)
  );
  GT_2x1 GT907 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1053:134
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup906__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1052:148
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1760_2700_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2718:150
    ._dfc_wire_2105                          (_GT907__dfc_wire_2105)
  );
  MUX_3x1 MUX908 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1054:163
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT907__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1053:134
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_27_2697_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2715:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1787_2698_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2716:150
    ._dfc_wire_2108                          (_MUX908__dfc_wire_2108)
  );
  LT_2x1 LT909 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1055:134
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup906__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1052:148
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1726_2696_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2714:150
    ._dfc_wire_2112                          (_LT909__dfc_wire_2112)
  );
  MUX_3x1 MUX910 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1056:163
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_36_2692_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2710:138
    ._dfc_wire_2103_2110                     (_MUX908__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1054:163
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1824_2693_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2711:150
    ._dfc_wire_2108                          (_MUX910__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST911 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1057:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX910__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1056:163
    ._dfc_wire_236 (sink__dfc_wire_2141__dfc_wire_4799)
  );
  dup_1x2 dup912 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1058:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB879__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1025:109
    ._dfc_wire_68_105 (_dup912__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup912__dfc_wire_68_113)
  );
  dup_1x2 dup913 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1059:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR8889__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1035:87
    ._dfc_wire_68_105 (_dup913__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup913__dfc_wire_68_113)
  );
  ADD_2x1 ADD914 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1060:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_342_2687_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2705:146
    .const_fix_32_0_1__0000000000000080_102 (_dup913__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1059:111
    ._dfc_wire_100                          (_ADD914__dfc_wire_100)
  );
  SHR14_1x1 SHR14915 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1061:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD914__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1060:130
    ._dfc_wire_2103 (_SHR14915__dfc_wire_2103)
  );
  dup_1x3 dup916 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1062:148
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR14915__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1061:93
    ._dfc_wire_2103_2106 (_dup916__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup916__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup916__dfc_wire_2103_2113)
  );
  GT_2x1 GT917 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1063:134
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup916__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1062:148
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1750_2684_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2702:150
    ._dfc_wire_2105                          (_GT917__dfc_wire_2105)
  );
  MUX_3x1 MUX918 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1064:163
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT917__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1063:134
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_19_2680_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2698:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1769_2681_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2699:150
    ._dfc_wire_2108                          (_MUX918__dfc_wire_2108)
  );
  LT_2x1 LT919 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1065:134
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup916__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1062:148
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1716_2678_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2696:150
    ._dfc_wire_2112                          (_LT919__dfc_wire_2112)
  );
  MUX_3x1 MUX920 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1066:163
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_27_2676_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2694:138
    ._dfc_wire_2103_2110                     (_MUX918__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1064:163
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1781_2677_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2695:150
    ._dfc_wire_2108                          (_MUX920__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST921 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1067:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX920__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1066:163
    ._dfc_wire_236 (sink__dfc_wire_2163__dfc_wire_4799)
  );
  dup_1x2 dup922 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1068:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB875__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1021:109
    ._dfc_wire_68_105 (_dup922__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup922__dfc_wire_68_113)
  );
  dup_1x2 dup923 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1069:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD870__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1016:130
    ._dfc_wire_68_105 (_dup923__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup923__dfc_wire_68_113)
  );
  ADD_2x1 ADD924 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1070:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_127_2669_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2687:146
    .const_fix_32_0_1__0000000000000080_102 (_dup923__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1069:111
    ._dfc_wire_100                          (_ADD924__dfc_wire_100)
  );
  SHR14_1x1 SHR14925 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1071:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD924__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1070:130
    ._dfc_wire_2103 (_SHR14925__dfc_wire_2103)
  );
  dup_1x3 dup926 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1072:148
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR14925__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1071:93
    ._dfc_wire_2103_2106 (_dup926__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup926__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup926__dfc_wire_2103_2113)
  );
  GT_2x1 GT927 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1073:134
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup926__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1072:148
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1433_2665_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2683:150
    ._dfc_wire_2105                          (_GT927__dfc_wire_2105)
  );
  MUX_3x1 MUX928 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1074:163
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT927__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1073:134
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_96_2661_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2679:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1529_2662_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2680:150
    ._dfc_wire_2108                          (_MUX928__dfc_wire_2108)
  );
  LT_2x1 LT929 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1075:134
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup926__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1072:148
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1399_2659_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2677:150
    ._dfc_wire_2112                          (_LT929__dfc_wire_2112)
  );
  MUX_3x1 MUX930 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1076:163
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_108_2656_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2674:142
    ._dfc_wire_2103_2110                     (_MUX928__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1074:163
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1550_2657_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2675:150
    ._dfc_wire_2108                          (_MUX930__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST931 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1077:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX930__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1076:163
    ._dfc_wire_236 (sink__dfc_wire_2185__dfc_wire_4799)
  );
  SUB_2x1 SUB932 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1078:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_127_2653_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2671:146
    ._dfc_wire_118    (_dup923__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1069:111
    ._dfc_wire_121    (_SUB932__dfc_wire_121)
  );
  SHR14_1x1 SHR14933 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1079:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB932__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1078:109
    ._dfc_wire_2103 (_SHR14933__dfc_wire_2103)
  );
  dup_1x3 dup934 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1080:148
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR14933__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1079:93
    ._dfc_wire_2103_2106 (_dup934__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup934__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup934__dfc_wire_2103_2113)
  );
  GT_2x1 GT935 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1081:134
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup934__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1080:148
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1545_2650_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2668:150
    ._dfc_wire_2105                          (_GT935__dfc_wire_2105)
  );
  MUX_3x1 MUX936 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1082:163
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT935__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1081:134
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_26_2647_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2665:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1571_2648_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2666:150
    ._dfc_wire_2108                          (_MUX936__dfc_wire_2108)
  );
  LT_2x1 LT937 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1083:134
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup934__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1080:148
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1511_2630_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2648:150
    ._dfc_wire_2112                          (_LT937__dfc_wire_2112)
  );
  MUX_3x1 MUX938 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1084:163
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_LT937__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1083:134
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_11_2628_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2646:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1575_2629_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2647:150
    ._dfc_wire_2108                          (_MUX938__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST939 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1085:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX938__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1084:163
    ._dfc_wire_236 (sink__dfc_wire_2207__dfc_wire_4799)
  );
  SUB_2x1 SUB940 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1086:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_342_2626_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2644:146
    ._dfc_wire_118    (_dup913__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1059:111
    ._dfc_wire_121    (_SUB940__dfc_wire_121)
  );
  SHR14_1x1 SHR14941 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1087:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB940__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1086:109
    ._dfc_wire_2103 (_SHR14941__dfc_wire_2103)
  );
  dup_1x3 dup942 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1088:148
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR14941__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1087:93
    ._dfc_wire_2103_2106 (_dup942__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup942__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup942__dfc_wire_2103_2113)
  );
  GT_2x1 GT943 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1089:134
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup942__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1088:148
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1736_2623_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2641:150
    ._dfc_wire_2105                          (_GT943__dfc_wire_2105)
  );
  MUX_3x1 MUX944 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1090:163
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT943__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1089:134
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_22_2620_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2638:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1758_2621_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2639:150
    ._dfc_wire_2108                          (_MUX944__dfc_wire_2108)
  );
  LT_2x1 LT945 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1091:134
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup942__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1088:148
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1702_2616_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2634:150
    ._dfc_wire_2112                          (_LT945__dfc_wire_2112)
  );
  MUX_3x1 MUX946 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1092:163
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_LT945__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1091:134
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_33_2613_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2631:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1758_2614_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2632:150
    ._dfc_wire_2108                          (_MUX946__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST947 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1093:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX946__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1092:163
    ._dfc_wire_236 (sink__dfc_wire_2229__dfc_wire_4799)
  );
  SUB_2x1 SUB948 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1094:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_460_2610_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2628:146
    ._dfc_wire_118    (_dup903__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1049:111
    ._dfc_wire_121    (_SUB948__dfc_wire_121)
  );
  SHR14_1x1 SHR14949 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1095:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB948__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1094:109
    ._dfc_wire_2103 (_SHR14949__dfc_wire_2103)
  );
  dup_1x3 dup950 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1096:148
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR14949__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1095:93
    ._dfc_wire_2103_2106 (_dup950__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup950__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup950__dfc_wire_2103_2113)
  );
  GT_2x1 GT951 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1097:134
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup950__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1096:148
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1915_2608_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2626:150
    ._dfc_wire_2105                          (_GT951__dfc_wire_2105)
  );
  MUX_3x1 MUX952 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1098:163
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT951__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1097:134
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_41_2606_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2624:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1956_2607_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2625:150
    ._dfc_wire_2108                          (_MUX952__dfc_wire_2108)
  );
  LT_2x1 LT953 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1099:134
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup950__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1096:148
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1881_2605_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2623:150
    ._dfc_wire_2112                          (_LT953__dfc_wire_2112)
  );
  MUX_3x1 MUX954 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1100:163
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_53_2602_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2620:138
    ._dfc_wire_2103_2110                     (_MUX952__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1098:163
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1963_2603_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2621:150
    ._dfc_wire_2108                          (_MUX954__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST955 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1101:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX954__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1100:163
    ._dfc_wire_236 (sink__dfc_wire_2251__dfc_wire_4799)
  );
  SUB_2x1 SUB956 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1102:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_190_2598_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2616:146
    ._dfc_wire_118    (_dup891__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1037:111
    ._dfc_wire_121    (_SUB956__dfc_wire_121)
  );
  SHR14_1x1 SHR14957 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1103:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB956__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1102:109
    ._dfc_wire_2103 (_SHR14957__dfc_wire_2103)
  );
  dup_1x3 dup958 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1104:148
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR14957__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1103:93
    ._dfc_wire_2103_2106 (_dup958__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup958__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup958__dfc_wire_2103_2113)
  );
  GT_2x1 GT959 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1105:134
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup958__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1104:148
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1604_2594_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2612:150
    ._dfc_wire_2105                          (_GT959__dfc_wire_2105)
  );
  MUX_3x1 MUX960 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1106:163
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT959__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1105:134
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_47_2592_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2610:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1651_2593_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2611:150
    ._dfc_wire_2108                          (_MUX960__dfc_wire_2108)
  );
  LT_2x1 LT961 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1107:134
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup958__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1104:148
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1570_2590_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2608:150
    ._dfc_wire_2112                          (_LT961__dfc_wire_2112)
  );
  MUX_3x1 MUX962 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1108:163
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_LT961__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1107:134
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_13_2587_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2605:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1666_2588_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2606:150
    ._dfc_wire_2108                          (_MUX962__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST963 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1109:87
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX962__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1108:163
    ._dfc_wire_236 (sink__dfc_wire_2273__dfc_wire_4799)
  );
  CAST_1x1_16_32 CAST964 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1110:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST488__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:634:87
    ._dfc_wire_73 (_CAST964__dfc_wire_73)
  );
  SHL8_1x1 SHL8965 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1111:89
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1921 (_CAST964__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1110:84
    ._dfc_wire_1923 (_SHL8965__dfc_wire_1923)
  );
  CAST_1x1_16_32 CAST966 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1112:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST688__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:834:87
    ._dfc_wire_73 (_CAST966__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST967 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1113:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST288__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:434:87
    ._dfc_wire_73 (_CAST967__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST968 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1114:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST188__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:334:87
    ._dfc_wire_73 (_CAST968__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST969 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1115:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST788__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:934:87
    ._dfc_wire_73 (_CAST969__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST970 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1116:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST588__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:734:87
    ._dfc_wire_73 (_CAST970__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST971 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1117:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST388__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:534:87
    ._dfc_wire_73 (_CAST971__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST972 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1118:84
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST88__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:234:83
    ._dfc_wire_73 (_CAST972__dfc_wire_73)
  );
  SHL8_1x1 SHL8973 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1119:89
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1921 (_CAST972__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1118:84
    ._dfc_wire_1923 (_SHL8973__dfc_wire_1923)
  );
  ADD_2x1 ADD974 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1120:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_SHL8973__dfc_wire_1923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1119:89
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1021_2574_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2592:150
    ._dfc_wire_100                          (_ADD974__dfc_wire_100)
  );
  dup_1x2 dup975 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1121:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST968__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1114:84
    ._dfc_wire_68_105 (_dup975__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup975__dfc_wire_68_113)
  );
  dup_1x2 dup976 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1122:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST969__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1115:84
    ._dfc_wire_68_105 (_dup976__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup976__dfc_wire_68_113)
  );
  ADD_2x1 ADD977 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1123:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup975__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1121:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_283_2566_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2584:146
    ._dfc_wire_100                          (_ADD977__dfc_wire_100)
  );
  MUL_2x1 MUL978 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1124:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1147_2564_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2582:150
    ._dfc_wire_104                          (_ADD977__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1123:130
    ._dfc_wire_107                          (_MUL978__dfc_wire_107)
  );
  ADD_2x1 ADD979 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1125:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL978__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1124:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1070_3066_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3084:150
    ._dfc_wire_100                          (_ADD979__dfc_wire_100)
  );
  MUL_2x1 MUL980 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1126:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1100_3065_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3083:150
    ._dfc_wire_104                          (_dup975__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1121:111
    ._dfc_wire_107                          (_MUL980__dfc_wire_107)
  );
  dup_1x2 dup981 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1127:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD979__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1125:130
    ._dfc_wire_68_105 (_dup981__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup981__dfc_wire_68_113)
  );
  ADD_2x1 ADD982 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1128:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup981__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1127:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_125_3060_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3078:146
    ._dfc_wire_100                          (_ADD982__dfc_wire_100)
  );
  SHR3_1x1 SHR3983 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1129:89
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_ADD982__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1128:130
    ._dfc_wire_1968 (_SHR3983__dfc_wire_1968)
  );
  MUL_2x1 MUL984 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1130:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_861_3054_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3072:146
    ._dfc_wire_104                          (_dup976__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1122:111
    ._dfc_wire_107                          (_MUL984__dfc_wire_107)
  );
  SUB_2x1 SUB985 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1131:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup981__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1127:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_386_3050_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3068:146
    ._dfc_wire_121    (_SUB985__dfc_wire_121)
  );
  SHR3_1x1 SHR3986 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1132:89
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB985__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1131:109
    ._dfc_wire_1968 (_SHR3986__dfc_wire_1968)
  );
  dup_1x2 dup987 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1133:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST970__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1116:84
    ._dfc_wire_68_105 (_dup987__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup987__dfc_wire_68_113)
  );
  dup_1x2 dup988 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1134:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST971__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1117:84
    ._dfc_wire_68_105 (_dup988__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup988__dfc_wire_68_113)
  );
  ADD_2x1 ADD989 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1135:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup987__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1133:111
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_87_3043_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3061:142
    ._dfc_wire_100                          (_ADD989__dfc_wire_100)
  );
  MUL_2x1 MUL990 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1136:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1099_3040_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3058:150
    ._dfc_wire_104                          (_ADD989__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1135:130
    ._dfc_wire_107                          (_MUL990__dfc_wire_107)
  );
  ADD_2x1 ADD991 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1137:130
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL990__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1136:131
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1076_3036_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3054:150
    ._dfc_wire_100                          (_ADD991__dfc_wire_100)
  );
  MUL_2x1 MUL992 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1138:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_983_3033_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3051:146
    ._dfc_wire_104                          (_dup987__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1133:111
    ._dfc_wire_107                          (_MUL992__dfc_wire_107)
  );
  dup_1x2 dup993 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1139:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD991__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1137:130
    ._dfc_wire_68_105 (_dup993__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup993__dfc_wire_68_113)
  );
  SUB_2x1 SUB994 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1140:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup993__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1139:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_246_3229_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3247:146
    ._dfc_wire_121    (_SUB994__dfc_wire_121)
  );
  SHR3_1x1 SHR3995 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1141:89
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB994__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1140:109
    ._dfc_wire_1968 (_SHR3995__dfc_wire_1968)
  );
  MUL_2x1 MUL996 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1142:131
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_954_3027_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3045:146
    ._dfc_wire_104                          (_dup988__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1134:111
    ._dfc_wire_107                          (_MUL996__dfc_wire_107)
  );
  SUB_2x1 SUB997 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1143:109
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup993__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1139:111
    ._dfc_wire_118    (_delay_fixed_32_0_1_359_3025_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3043:146
    ._dfc_wire_121    (_SUB997__dfc_wire_121)
  );
  SHR3_1x1 SHR3998 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1144:89
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB997__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1143:109
    ._dfc_wire_1968 (_SHR3998__dfc_wire_1968)
  );
  dup_1x2 dup999 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1145:111
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD974__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1120:130
    ._dfc_wire_68_105 (_dup999__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup999__dfc_wire_68_113)
  );
  dup_1x2 dup1000 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1146:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHL8965__dfc_wire_1923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1111:89
    ._dfc_wire_68_105 (_dup1000__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1000__dfc_wire_68_113)
  );
  ADD_2x1 ADD1001 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1147:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_25_3015_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3033:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1000__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1146:116
    ._dfc_wire_100                          (_ADD1001__dfc_wire_100)
  );
  SUB_2x1 SUB1002 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1148:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_25_3014_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3032:142
    ._dfc_wire_118    (_dup1000__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1146:116
    ._dfc_wire_121    (_SUB1002__dfc_wire_121)
  );
  dup_1x2 dup1003 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1149:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST967__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1113:84
    ._dfc_wire_68_105 (_dup1003__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1003__dfc_wire_68_113)
  );
  dup_1x2 dup1004 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1150:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST966__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1112:84
    ._dfc_wire_68_105 (_dup1004__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1004__dfc_wire_68_113)
  );
  ADD_2x1 ADD1005 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1151:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1003__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1149:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_287_3009_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3027:146
    ._dfc_wire_100                          (_ADD1005__dfc_wire_100)
  );
  MUL_2x1 MUL1006 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1152:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1037_3007_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3025:150
    ._dfc_wire_104                          (_ADD1005__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1151:135
    ._dfc_wire_107                          (_MUL1006__dfc_wire_107)
  );
  ADD_2x1 ADD1007 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1153:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1006__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1152:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_966_3004_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3022:146
    ._dfc_wire_100                          (_ADD1007__dfc_wire_100)
  );
  MUL_2x1 MUL1008 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1154:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_689_3001_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3019:146
    ._dfc_wire_104                          (_dup1004__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1150:116
    ._dfc_wire_107                          (_MUL1008__dfc_wire_107)
  );
  dup_1x2 dup1009 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1155:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1007__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1153:135
    ._dfc_wire_68_105 (_dup1009__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1009__dfc_wire_68_113)
  );
  SUB_2x1 SUB1010 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1156:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1009__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1155:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_461_2996_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3014:146
    ._dfc_wire_121    (_SUB1010__dfc_wire_121)
  );
  SHR3_1x1 SHR31011 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1157:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1010__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1156:114
    ._dfc_wire_1968 (_SHR31011__dfc_wire_1968)
  );
  MUL_2x1 MUL1012 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1158:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1032_2994_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3012:150
    ._dfc_wire_104                          (_dup1003__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1149:116
    ._dfc_wire_107                          (_MUL1012__dfc_wire_107)
  );
  ADD_2x1 ADD1013 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1159:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1009__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1155:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_128_3210_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3228:146
    ._dfc_wire_100                          (_ADD1013__dfc_wire_100)
  );
  SHR3_1x1 SHR31014 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1160:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_ADD1013__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1159:135
    ._dfc_wire_1968 (_SHR31014__dfc_wire_1968)
  );
  dup_1x2 dup1015 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1161:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR3983__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1129:89
    ._dfc_wire_68_105 (_dup1015__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1015__dfc_wire_68_113)
  );
  dup_1x2 dup1016 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1162:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR3995__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1141:89
    ._dfc_wire_68_105 (_dup1016__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1016__dfc_wire_68_113)
  );
  ADD_2x1 ADD1017 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1163:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1015__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1161:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_4_2990_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3008:138
    ._dfc_wire_100                          (_ADD1017__dfc_wire_100)
  );
  SUB_2x1 SUB1018 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1164:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1015__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1161:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_4_2989_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3007:138
    ._dfc_wire_121    (_SUB1018__dfc_wire_121)
  );
  dup_1x2 dup1019 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1165:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR3986__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1132:89
    ._dfc_wire_68_105 (_dup1019__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1019__dfc_wire_68_113)
  );
  dup_1x2 dup1020 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1166:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR3998__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1144:89
    ._dfc_wire_68_105 (_dup1020__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1020__dfc_wire_68_113)
  );
  ADD_2x1 ADD1021 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1167:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_70_2985_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3003:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1020__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1166:116
    ._dfc_wire_100                          (_ADD1021__dfc_wire_100)
  );
  SUB_2x1 SUB1022 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1168:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_70_2982_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3000:142
    ._dfc_wire_118    (_dup1020__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1166:116
    ._dfc_wire_121    (_SUB1022__dfc_wire_121)
  );
  dup_1x2 dup1023 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1169:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1001__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1147:135
    ._dfc_wire_68_105 (_dup1023__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1023__dfc_wire_68_113)
  );
  dup_1x2 dup1024 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1170:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31014__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1160:93
    ._dfc_wire_68_105 (_dup1024__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1024__dfc_wire_68_113)
  );
  ADD_2x1 ADD1025 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1171:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_256_2560_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2578:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1024__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1170:116
    ._dfc_wire_100                          (_ADD1025__dfc_wire_100)
  );
  SUB_2x1 SUB1026 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1172:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_256_2559_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2577:146
    ._dfc_wire_118    (_dup1024__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1170:116
    ._dfc_wire_121    (_SUB1026__dfc_wire_121)
  );
  dup_1x2 dup1027 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1173:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1002__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1148:114
    ._dfc_wire_68_105 (_dup1027__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1027__dfc_wire_68_113)
  );
  dup_1x2 dup1028 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1174:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31011__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1157:93
    ._dfc_wire_68_105 (_dup1028__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1028__dfc_wire_68_113)
  );
  ADD_2x1 ADD1029 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1175:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_226_2558_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2576:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1028__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1174:116
    ._dfc_wire_100                          (_ADD1029__dfc_wire_100)
  );
  SUB_2x1 SUB1030 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1176:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_226_2557_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2575:146
    ._dfc_wire_118    (_dup1028__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1174:116
    ._dfc_wire_121    (_SUB1030__dfc_wire_121)
  );
  dup_1x2 dup1031 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1177:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1018__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1164:114
    ._dfc_wire_68_105 (_dup1031__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1031__dfc_wire_68_113)
  );
  dup_1x2 dup1032 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1178:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1022__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1168:114
    ._dfc_wire_68_105 (_dup1032__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1032__dfc_wire_68_113)
  );
  ADD_2x1 ADD1033 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1179:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1031__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1177:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_80_2556_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2574:142
    ._dfc_wire_100                          (_ADD1033__dfc_wire_100)
  );
  MUL_2x1 MUL1034 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1180:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1728_2555_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2573:150
    ._dfc_wire_104                          (_ADD1033__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1179:135
    ._dfc_wire_107                          (_MUL1034__dfc_wire_107)
  );
  ADD_2x1 ADD1035 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1181:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1034__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1180:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1838_2554_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2572:150
    ._dfc_wire_100                          (_ADD1035__dfc_wire_100)
  );
  SHR8_1x1 SHR81036 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1182:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD1035__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1181:135
    ._dfc_wire_216 (_SHR81036__dfc_wire_216)
  );
  SUB_2x1 SUB1037 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1183:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1031__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1177:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_80_2553_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2571:142
    ._dfc_wire_121    (_SUB1037__dfc_wire_121)
  );
  MUL_2x1 MUL1038 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1184:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1732_2552_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2570:150
    ._dfc_wire_104                          (_SUB1037__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1183:114
    ._dfc_wire_107                          (_MUL1038__dfc_wire_107)
  );
  ADD_2x1 ADD1039 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1185:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1038__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1184:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1811_2551_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2569:150
    ._dfc_wire_100                          (_ADD1039__dfc_wire_100)
  );
  SHR8_1x1 SHR81040 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1186:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD1039__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1185:135
    ._dfc_wire_216 (_SHR81040__dfc_wire_216)
  );
  dup_1x2 dup1041 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1187:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1025__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1171:135
    ._dfc_wire_68_105 (_dup1041__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1041__dfc_wire_68_113)
  );
  dup_1x2 dup1042 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1188:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1017__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1163:135
    ._dfc_wire_68_105 (_dup1042__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1042__dfc_wire_68_113)
  );
  ADD_2x1 ADD1043 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1189:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_59_2550_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2568:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1042__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1188:116
    ._dfc_wire_100                          (_ADD1043__dfc_wire_100)
  );
  SHR14_1x1 SHR141044 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1190:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1043__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1189:135
    ._dfc_wire_2103 (_SHR141044__dfc_wire_2103)
  );
  dup_1x3 dup1045 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1191:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141044__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1190:97
    ._dfc_wire_2103_2106 (_dup1045__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1045__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1045__dfc_wire_2103_2113)
  );
  GT_2x1 GT1046 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1192:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1045__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1191:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1747_2549_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2567:150
    ._dfc_wire_2105                          (_GT1046__dfc_wire_2105)
  );
  MUX_3x1 MUX1047 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1193:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1046__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1192:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_39_2547_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2565:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1786_2548_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2566:150
    ._dfc_wire_2108                          (_MUX1047__dfc_wire_2108)
  );
  LT_2x1 LT1048 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1194:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1045__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1191:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1713_2546_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2564:150
    ._dfc_wire_2112                          (_LT1048__dfc_wire_2112)
  );
  MUX_3x1 MUX1049 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1195:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_75_2544_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2562:138
    ._dfc_wire_2103_2110                     (_MUX1047__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1193:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1807_2545_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2563:150
    ._dfc_wire_2108                          (_MUX1049__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1050 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1196:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1049__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1195:169
    ._dfc_wire_236 (sink__dfc_wire_2483__dfc_wire_4799)
  );
  dup_1x2 dup1051 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1197:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1029__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1175:135
    ._dfc_wire_68_105 (_dup1051__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1051__dfc_wire_68_113)
  );
  dup_1x2 dup1052 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1198:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR81036__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1182:91
    ._dfc_wire_68_105 (_dup1052__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1052__dfc_wire_68_113)
  );
  ADD_2x1 ADD1053 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1199:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_478_2543_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2561:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1052__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1198:116
    ._dfc_wire_100                          (_ADD1053__dfc_wire_100)
  );
  SHR14_1x1 SHR141054 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1200:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1053__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1199:135
    ._dfc_wire_2103 (_SHR141054__dfc_wire_2103)
  );
  dup_1x3 dup1055 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1201:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141054__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1200:97
    ._dfc_wire_2103_2106 (_dup1055__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1055__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1055__dfc_wire_2103_2113)
  );
  GT_2x1 GT1056 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1202:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1055__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1201:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_2173_2542_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2560:150
    ._dfc_wire_2105                          (_GT1056__dfc_wire_2105)
  );
  MUX_3x1 MUX1057 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1203:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1056__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1202:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_89_2540_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2558:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_2262_2541_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2559:150
    ._dfc_wire_2108                          (_MUX1057__dfc_wire_2108)
  );
  LT_2x1 LT1058 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1204:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1055__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1201:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_2139_2539_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2557:150
    ._dfc_wire_2112                          (_LT1058__dfc_wire_2112)
  );
  MUX_3x1 MUX1059 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1205:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_85_3175_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3193:138
    ._dfc_wire_2103_2110                     (_MUX1057__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1203:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_2274_3176_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3194:150
    ._dfc_wire_2108                          (_MUX1059__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1060 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1206:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1059__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1205:169
    ._dfc_wire_236 (sink__dfc_wire_2505__dfc_wire_4799)
  );
  dup_1x2 dup1061 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1207:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1030__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1176:114
    ._dfc_wire_68_105 (_dup1061__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1061__dfc_wire_68_113)
  );
  dup_1x2 dup1062 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1208:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR81040__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1186:91
    ._dfc_wire_68_105 (_dup1062__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1062__dfc_wire_68_113)
  );
  ADD_2x1 ADD1063 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1209:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_365_3173_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3191:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1062__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1208:116
    ._dfc_wire_100                          (_ADD1063__dfc_wire_100)
  );
  SHR14_1x1 SHR141064 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1210:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1063__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1209:135
    ._dfc_wire_2103 (_SHR141064__dfc_wire_2103)
  );
  dup_1x3 dup1065 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1211:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141064__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1210:97
    ._dfc_wire_2103_2106 (_dup1065__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1065__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1065__dfc_wire_2103_2113)
  );
  GT_2x1 GT1066 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1212:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1065__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1211:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1987_3171_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3189:150
    ._dfc_wire_2105                          (_GT1066__dfc_wire_2105)
  );
  MUX_3x1 MUX1067 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1213:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1066__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1212:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_4_3168_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3186:138
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1991_3169_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3187:150
    ._dfc_wire_2108                          (_MUX1067__dfc_wire_2108)
  );
  LT_2x1 LT1068 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1214:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1065__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1211:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1953_3167_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3185:150
    ._dfc_wire_2112                          (_LT1068__dfc_wire_2112)
  );
  MUX_3x1 MUX1069 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1215:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_2_3165_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3183:134
    ._dfc_wire_2103_2110                     (_MUX1067__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1213:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_2006_3166_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3184:150
    ._dfc_wire_2108                          (_MUX1069__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1070 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1216:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1069__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1215:169
    ._dfc_wire_236 (sink__dfc_wire_2527__dfc_wire_4799)
  );
  dup_1x2 dup1071 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1217:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1026__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1172:114
    ._dfc_wire_68_105 (_dup1071__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1071__dfc_wire_68_113)
  );
  dup_1x2 dup1072 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1218:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1021__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1167:135
    ._dfc_wire_68_105 (_dup1072__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1072__dfc_wire_68_113)
  );
  ADD_2x1 ADD1073 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1219:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_156_3164_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3182:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1072__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1218:116
    ._dfc_wire_100                          (_ADD1073__dfc_wire_100)
  );
  SHR14_1x1 SHR141074 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1220:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1073__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1219:135
    ._dfc_wire_2103 (_SHR141074__dfc_wire_2103)
  );
  dup_1x3 dup1075 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1221:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141074__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1220:97
    ._dfc_wire_2103_2106 (_dup1075__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1075__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1075__dfc_wire_2103_2113)
  );
  GT_2x1 GT1076 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1222:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1075__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1221:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1796_3163_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3181:150
    ._dfc_wire_2105                          (_GT1076__dfc_wire_2105)
  );
  MUX_3x1 MUX1077 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1223:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1076__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1222:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_39_3161_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3179:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1835_3162_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3180:150
    ._dfc_wire_2108                          (_MUX1077__dfc_wire_2108)
  );
  LT_2x1 LT1078 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1224:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1075__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1221:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1762_3160_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3178:150
    ._dfc_wire_2112                          (_LT1078__dfc_wire_2112)
  );
  MUX_3x1 MUX1079 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1225:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_52_3158_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3176:138
    ._dfc_wire_2103_2110                     (_MUX1077__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1223:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1895_3159_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3177:150
    ._dfc_wire_2108                          (_MUX1079__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1080 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1226:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1079__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1225:169
    ._dfc_wire_236 (sink__dfc_wire_2549__dfc_wire_4799)
  );
  SUB_2x1 SUB1081 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1227:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_156_3156_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3174:146
    ._dfc_wire_118    (_dup1072__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1218:116
    ._dfc_wire_121    (_SUB1081__dfc_wire_121)
  );
  SHR14_1x1 SHR141082 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1228:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1081__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1227:114
    ._dfc_wire_2103 (_SHR141082__dfc_wire_2103)
  );
  dup_1x3 dup1083 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1229:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141082__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1228:97
    ._dfc_wire_2103_2106 (_dup1083__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1083__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1083__dfc_wire_2103_2113)
  );
  GT_2x1 GT1084 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1230:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1083__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1229:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1713_3153_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3171:150
    ._dfc_wire_2105                          (_GT1084__dfc_wire_2105)
  );
  MUX_3x1 MUX1085 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1231:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1084__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1230:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_71_3150_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3168:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1784_3151_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3169:150
    ._dfc_wire_2108                          (_MUX1085__dfc_wire_2108)
  );
  LT_2x1 LT1086 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1232:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1083__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1229:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1679_3149_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3167:150
    ._dfc_wire_2112                          (_LT1086__dfc_wire_2112)
  );
  MUX_3x1 MUX1087 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1233:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_30_3146_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3164:138
    ._dfc_wire_2103_2110                     (_MUX1085__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1231:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1774_3147_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3165:150
    ._dfc_wire_2108                          (_MUX1087__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1088 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1234:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1087__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1233:169
    ._dfc_wire_236 (sink__dfc_wire_2571__dfc_wire_4799)
  );
  SUB_2x1 SUB1089 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1235:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_365_3078_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3096:146
    ._dfc_wire_118    (_dup1062__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1208:116
    ._dfc_wire_121    (_SUB1089__dfc_wire_121)
  );
  SHR14_1x1 SHR141090 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1236:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1089__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1235:114
    ._dfc_wire_2103 (_SHR141090__dfc_wire_2103)
  );
  dup_1x3 dup1091 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1237:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141090__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1236:97
    ._dfc_wire_2103_2106 (_dup1091__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1091__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1091__dfc_wire_2103_2113)
  );
  GT_2x1 GT1092 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1238:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1091__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1237:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_2076_3075_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3093:150
    ._dfc_wire_2105                          (_GT1092__dfc_wire_2105)
  );
  MUX_3x1 MUX1093 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1239:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1092__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1238:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_63_3073_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3091:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_2139_3074_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3092:150
    ._dfc_wire_2108                          (_MUX1093__dfc_wire_2108)
  );
  LT_2x1 LT1094 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1240:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1091__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1237:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_2042_3071_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3089:150
    ._dfc_wire_2112                          (_LT1094__dfc_wire_2112)
  );
  MUX_3x1 MUX1095 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1241:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_60_3068_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3086:138
    ._dfc_wire_2103_2110                     (_MUX1093__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1239:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_2172_3069_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3087:150
    ._dfc_wire_2108                          (_MUX1095__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1096 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1242:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1095__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1241:169
    ._dfc_wire_236 (sink__dfc_wire_2593__dfc_wire_4799)
  );
  SUB_2x1 SUB1097 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1243:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_478_2538_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2556:146
    ._dfc_wire_118    (_dup1052__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1198:116
    ._dfc_wire_121    (_SUB1097__dfc_wire_121)
  );
  SHR14_1x1 SHR141098 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1244:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1097__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1243:114
    ._dfc_wire_2103 (_SHR141098__dfc_wire_2103)
  );
  dup_1x3 dup1099 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1245:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141098__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1244:97
    ._dfc_wire_2103_2106 (_dup1099__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1099__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1099__dfc_wire_2103_2113)
  );
  GT_2x1 GT1100 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1246:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1099__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1245:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_2078_2537_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2555:150
    ._dfc_wire_2105                          (_GT1100__dfc_wire_2105)
  );
  MUX_3x1 MUX1101 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1247:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1100__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1246:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_7_2535_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2553:138
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_2085_2536_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2554:150
    ._dfc_wire_2108                          (_MUX1101__dfc_wire_2108)
  );
  LT_2x1 LT1102 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1248:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1099__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1245:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_2044_2534_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2552:150
    ._dfc_wire_2112                          (_LT1102__dfc_wire_2112)
  );
  MUX_3x1 MUX1103 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1249:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_9_2532_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2550:134
    ._dfc_wire_2103_2110                     (_MUX1101__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1247:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_2086_2533_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2551:150
    ._dfc_wire_2108                          (_MUX1103__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1104 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1250:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1103__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1249:169
    ._dfc_wire_236 (sink__dfc_wire_2615__dfc_wire_4799)
  );
  SUB_2x1 SUB1105 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1251:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_59_2531_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2549:142
    ._dfc_wire_118    (_dup1042__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1188:116
    ._dfc_wire_121    (_SUB1105__dfc_wire_121)
  );
  SHR14_1x1 SHR141106 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1252:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1105__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1251:114
    ._dfc_wire_2103 (_SHR141106__dfc_wire_2103)
  );
  dup_1x3 dup1107 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1253:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141106__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1252:97
    ._dfc_wire_2103_2106 (_dup1107__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1107__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1107__dfc_wire_2103_2113)
  );
  GT_2x1 GT1108 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1254:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1107__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1253:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1678_2530_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2548:150
    ._dfc_wire_2105                          (_GT1108__dfc_wire_2105)
  );
  MUX_3x1 MUX1109 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1255:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1108__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1254:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_39_2528_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2546:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1717_2529_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2547:150
    ._dfc_wire_2108                          (_MUX1109__dfc_wire_2108)
  );
  LT_2x1 LT1110 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1256:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1107__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1253:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1644_2527_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2545:150
    ._dfc_wire_2112                          (_LT1110__dfc_wire_2112)
  );
  MUX_3x1 MUX1111 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1257:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_95_2525_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2543:138
    ._dfc_wire_2103_2110                     (_MUX1109__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1255:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1777_2526_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2544:150
    ._dfc_wire_2108                          (_MUX1111__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1112 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1258:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1111__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1257:169
    ._dfc_wire_236 (sink__dfc_wire_2637__dfc_wire_4799)
  );
  CAST_1x1_16_32 CAST1113 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1259:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST493__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:639:87
    ._dfc_wire_73 (_CAST1113__dfc_wire_73)
  );
  SHL8_1x1 SHL81114 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1260:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1921 (_CAST1113__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1259:88
    ._dfc_wire_1923 (_SHL81114__dfc_wire_1923)
  );
  CAST_1x1_16_32 CAST1115 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1261:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST693__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:839:87
    ._dfc_wire_73 (_CAST1115__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1116 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1262:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST293__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:439:87
    ._dfc_wire_73 (_CAST1116__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1117 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1263:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST193__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:339:87
    ._dfc_wire_73 (_CAST1117__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1118 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1264:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST793__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:939:87
    ._dfc_wire_73 (_CAST1118__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1119 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1265:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST593__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:739:87
    ._dfc_wire_73 (_CAST1119__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1120 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1266:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST393__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:539:87
    ._dfc_wire_73 (_CAST1120__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1121 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1267:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST93__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:239:83
    ._dfc_wire_73 (_CAST1121__dfc_wire_73)
  );
  SHL8_1x1 SHL81122 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1268:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1921 (_CAST1121__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1267:88
    ._dfc_wire_1923 (_SHL81122__dfc_wire_1923)
  );
  ADD_2x1 ADD1123 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1269:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_SHL81122__dfc_wire_1923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1268:93
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_915_2524_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2542:146
    ._dfc_wire_100                          (_ADD1123__dfc_wire_100)
  );
  dup_1x2 dup1124 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1270:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1117__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1263:88
    ._dfc_wire_68_105 (_dup1124__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1124__dfc_wire_68_113)
  );
  dup_1x2 dup1125 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1271:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1118__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1264:88
    ._dfc_wire_68_105 (_dup1125__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1125__dfc_wire_68_113)
  );
  ADD_2x1 ADD1126 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1272:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_155_2523_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2541:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1125__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1271:116
    ._dfc_wire_100                          (_ADD1126__dfc_wire_100)
  );
  MUL_2x1 MUL1127 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1273:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1014_2522_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2540:150
    ._dfc_wire_104                          (_ADD1126__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1272:135
    ._dfc_wire_107                          (_MUL1127__dfc_wire_107)
  );
  ADD_2x1 ADD1128 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1274:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1127__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1273:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_983_2521_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2539:146
    ._dfc_wire_100                          (_ADD1128__dfc_wire_100)
  );
  MUL_2x1 MUL1129 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1275:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_781_2520_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2538:146
    ._dfc_wire_104                          (_dup1124__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1270:116
    ._dfc_wire_107                          (_MUL1129__dfc_wire_107)
  );
  dup_1x2 dup1130 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1276:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1128__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1274:135
    ._dfc_wire_68_105 (_dup1130__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1130__dfc_wire_68_113)
  );
  ADD_2x1 ADD1131 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1277:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1130__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1276:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_295_2519_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2537:146
    ._dfc_wire_100                          (_ADD1131__dfc_wire_100)
  );
  SHR3_1x1 SHR31132 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1278:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_ADD1131__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1277:135
    ._dfc_wire_1968 (_SHR31132__dfc_wire_1968)
  );
  MUL_2x1 MUL1133 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1279:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_980_2518_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2536:146
    ._dfc_wire_104                          (_dup1125__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1271:116
    ._dfc_wire_107                          (_MUL1133__dfc_wire_107)
  );
  SUB_2x1 SUB1134 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1280:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1130__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1276:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_138_2517_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2535:146
    ._dfc_wire_121    (_SUB1134__dfc_wire_121)
  );
  SHR3_1x1 SHR31135 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1281:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1134__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1280:114
    ._dfc_wire_1968 (_SHR31135__dfc_wire_1968)
  );
  dup_1x2 dup1136 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1282:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1119__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1265:88
    ._dfc_wire_68_105 (_dup1136__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1136__dfc_wire_68_113)
  );
  dup_1x2 dup1137 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1283:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1120__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1266:88
    ._dfc_wire_68_105 (_dup1137__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1137__dfc_wire_68_113)
  );
  ADD_2x1 ADD1138 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1284:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1136__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1282:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_73_2516_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2534:142
    ._dfc_wire_100                          (_ADD1138__dfc_wire_100)
  );
  MUL_2x1 MUL1139 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1285:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1032_2515_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2533:150
    ._dfc_wire_104                          (_ADD1138__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1284:135
    ._dfc_wire_107                          (_MUL1139__dfc_wire_107)
  );
  ADD_2x1 ADD1140 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1286:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1139__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1285:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1009_2514_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2532:150
    ._dfc_wire_100                          (_ADD1140__dfc_wire_100)
  );
  MUL_2x1 MUL1141 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1287:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_920_2513_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2531:146
    ._dfc_wire_104                          (_dup1136__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1282:116
    ._dfc_wire_107                          (_MUL1141__dfc_wire_107)
  );
  dup_1x2 dup1142 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1288:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1140__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1286:135
    ._dfc_wire_68_105 (_dup1142__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1142__dfc_wire_68_113)
  );
  SUB_2x1 SUB1143 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1289:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1142__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1288:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_222_3206_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3224:146
    ._dfc_wire_121    (_SUB1143__dfc_wire_121)
  );
  SHR3_1x1 SHR31144 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1290:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1143__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1289:114
    ._dfc_wire_1968 (_SHR31144__dfc_wire_1968)
  );
  MUL_2x1 MUL1145 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1291:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_905_3203_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3221:146
    ._dfc_wire_104                          (_dup1137__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1283:116
    ._dfc_wire_107                          (_MUL1145__dfc_wire_107)
  );
  SUB_2x1 SUB1146 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1292:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1142__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1288:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_259_3202_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3220:146
    ._dfc_wire_121    (_SUB1146__dfc_wire_121)
  );
  SHR3_1x1 SHR31147 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1293:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1146__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1292:114
    ._dfc_wire_1968 (_SHR31147__dfc_wire_1968)
  );
  dup_1x2 dup1148 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1294:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1123__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1269:135
    ._dfc_wire_68_105 (_dup1148__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1148__dfc_wire_68_113)
  );
  dup_1x2 dup1149 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1295:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHL81114__dfc_wire_1923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1260:93
    ._dfc_wire_68_105 (_dup1149__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1149__dfc_wire_68_113)
  );
  ADD_2x1 ADD1150 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1296:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1148__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1294:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_122_3106_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3124:146
    ._dfc_wire_100                          (_ADD1150__dfc_wire_100)
  );
  SUB_2x1 SUB1151 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1297:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1148__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1294:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_122_2512_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2530:146
    ._dfc_wire_121    (_SUB1151__dfc_wire_121)
  );
  dup_1x2 dup1152 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1298:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1116__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1262:88
    ._dfc_wire_68_105 (_dup1152__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1152__dfc_wire_68_113)
  );
  dup_1x2 dup1153 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1299:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1115__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1261:88
    ._dfc_wire_68_105 (_dup1153__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1153__dfc_wire_68_113)
  );
  ADD_2x1 ADD1154 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1300:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_7_2511_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2529:138
    .const_fix_32_0_1__0000000000000080_102 (_dup1153__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1299:116
    ._dfc_wire_100                          (_ADD1154__dfc_wire_100)
  );
  MUL_2x1 MUL1155 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1301:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1062_2510_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2528:150
    ._dfc_wire_104                          (_ADD1154__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1300:135
    ._dfc_wire_107                          (_MUL1155__dfc_wire_107)
  );
  ADD_2x1 ADD1156 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1302:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1155__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1301:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_986_2509_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2527:146
    ._dfc_wire_100                          (_ADD1156__dfc_wire_100)
  );
  MUL_2x1 MUL1157 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1303:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_994_2508_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2526:146
    ._dfc_wire_104                          (_dup1153__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1299:116
    ._dfc_wire_107                          (_MUL1157__dfc_wire_107)
  );
  dup_1x2 dup1158 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1304:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1156__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1302:135
    ._dfc_wire_68_105 (_dup1158__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1158__dfc_wire_68_113)
  );
  SUB_2x1 SUB1159 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1305:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1158__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1304:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_123_2507_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2525:146
    ._dfc_wire_121    (_SUB1159__dfc_wire_121)
  );
  SHR3_1x1 SHR31160 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1306:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1159__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1305:114
    ._dfc_wire_1968 (_SHR31160__dfc_wire_1968)
  );
  MUL_2x1 MUL1161 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1307:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1043_2506_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2524:150
    ._dfc_wire_104                          (_dup1152__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1298:116
    ._dfc_wire_107                          (_MUL1161__dfc_wire_107)
  );
  ADD_2x1 ADD1162 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1308:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1158__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1304:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_167_2505_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2523:146
    ._dfc_wire_100                          (_ADD1162__dfc_wire_100)
  );
  SHR3_1x1 SHR31163 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1309:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_ADD1162__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1308:135
    ._dfc_wire_1968 (_SHR31163__dfc_wire_1968)
  );
  dup_1x2 dup1164 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1310:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31132__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1278:93
    ._dfc_wire_68_105 (_dup1164__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1164__dfc_wire_68_113)
  );
  dup_1x2 dup1165 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1311:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31144__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1290:93
    ._dfc_wire_68_105 (_dup1165__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1165__dfc_wire_68_113)
  );
  ADD_2x1 ADD1166 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1312:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1164__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1310:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1_2504_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2522:138
    ._dfc_wire_100                          (_ADD1166__dfc_wire_100)
  );
  SUB_2x1 SUB1167 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1313:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1164__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1310:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_1_2503_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2521:138
    ._dfc_wire_121    (_SUB1167__dfc_wire_121)
  );
  dup_1x2 dup1168 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1314:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31135__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1281:93
    ._dfc_wire_68_105 (_dup1168__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1168__dfc_wire_68_113)
  );
  dup_1x2 dup1169 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1315:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31147__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1293:93
    ._dfc_wire_68_105 (_dup1169__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1169__dfc_wire_68_113)
  );
  ADD_2x1 ADD1170 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1316:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_25_2502_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2520:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1169__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1315:116
    ._dfc_wire_100                          (_ADD1170__dfc_wire_100)
  );
  SUB_2x1 SUB1171 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1317:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_25_2501_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2519:142
    ._dfc_wire_118    (_dup1169__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1315:116
    ._dfc_wire_121    (_SUB1171__dfc_wire_121)
  );
  dup_1x2 dup1172 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1318:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1150__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1296:135
    ._dfc_wire_68_105 (_dup1172__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1172__dfc_wire_68_113)
  );
  dup_1x2 dup1173 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1319:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31163__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1309:93
    ._dfc_wire_68_105 (_dup1173__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1173__dfc_wire_68_113)
  );
  ADD_2x1 ADD1174 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1320:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_270_2500_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2518:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1173__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1319:116
    ._dfc_wire_100                          (_ADD1174__dfc_wire_100)
  );
  SUB_2x1 SUB1175 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1321:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_270_2499_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2517:146
    ._dfc_wire_118    (_dup1173__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1319:116
    ._dfc_wire_121    (_SUB1175__dfc_wire_121)
  );
  dup_1x2 dup1176 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1322:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1151__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1297:114
    ._dfc_wire_68_105 (_dup1176__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1176__dfc_wire_68_113)
  );
  dup_1x2 dup1177 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1323:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31160__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1306:93
    ._dfc_wire_68_105 (_dup1177__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1177__dfc_wire_68_113)
  );
  ADD_2x1 ADD1178 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1324:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_172_2498_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2516:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1177__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1323:116
    ._dfc_wire_100                          (_ADD1178__dfc_wire_100)
  );
  SUB_2x1 SUB1179 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1325:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_172_2497_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2515:146
    ._dfc_wire_118    (_dup1177__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1323:116
    ._dfc_wire_121    (_SUB1179__dfc_wire_121)
  );
  dup_1x2 dup1180 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1326:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1167__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1313:114
    ._dfc_wire_68_105 (_dup1180__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1180__dfc_wire_68_113)
  );
  dup_1x2 dup1181 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1327:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1171__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1317:114
    ._dfc_wire_68_105 (_dup1181__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1181__dfc_wire_68_113)
  );
  ADD_2x1 ADD1182 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1328:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1180__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1326:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_111_2496_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2514:146
    ._dfc_wire_100                          (_ADD1182__dfc_wire_100)
  );
  MUL_2x1 MUL1183 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1329:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1578_2495_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2513:150
    ._dfc_wire_104                          (_ADD1182__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1328:135
    ._dfc_wire_107                          (_MUL1183__dfc_wire_107)
  );
  ADD_2x1 ADD1184 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1330:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1183__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1329:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1687_2494_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2512:150
    ._dfc_wire_100                          (_ADD1184__dfc_wire_100)
  );
  SHR8_1x1 SHR81185 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1331:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD1184__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1330:135
    ._dfc_wire_216 (_SHR81185__dfc_wire_216)
  );
  SUB_2x1 SUB1186 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1332:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1180__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1326:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_111_2493_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2511:146
    ._dfc_wire_121    (_SUB1186__dfc_wire_121)
  );
  MUL_2x1 MUL1187 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1333:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1556_2492_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2510:150
    ._dfc_wire_104                          (_SUB1186__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1332:114
    ._dfc_wire_107                          (_MUL1187__dfc_wire_107)
  );
  ADD_2x1 ADD1188 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1334:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1187__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1333:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1679_2491_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2509:150
    ._dfc_wire_100                          (_ADD1188__dfc_wire_100)
  );
  SHR8_1x1 SHR81189 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1335:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD1188__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1334:135
    ._dfc_wire_216 (_SHR81189__dfc_wire_216)
  );
  dup_1x2 dup1190 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1336:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1174__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1320:135
    ._dfc_wire_68_105 (_dup1190__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1190__dfc_wire_68_113)
  );
  dup_1x2 dup1191 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1337:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1166__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1312:135
    ._dfc_wire_68_105 (_dup1191__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1191__dfc_wire_68_113)
  );
  ADD_2x1 ADD1192 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1338:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_102_2490_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2508:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1191__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1337:116
    ._dfc_wire_100                          (_ADD1192__dfc_wire_100)
  );
  SHR14_1x1 SHR141193 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1339:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1192__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1338:135
    ._dfc_wire_2103 (_SHR141193__dfc_wire_2103)
  );
  dup_1x3 dup1194 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1340:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141193__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1339:97
    ._dfc_wire_2103_2106 (_dup1194__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1194__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1194__dfc_wire_2103_2113)
  );
  GT_2x1 GT1195 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1341:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1194__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1340:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1726_2489_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2507:150
    ._dfc_wire_2105                          (_GT1195__dfc_wire_2105)
  );
  MUX_3x1 MUX1196 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1342:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1195__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1341:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_92_2487_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2505:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1818_2488_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2506:150
    ._dfc_wire_2108                          (_MUX1196__dfc_wire_2108)
  );
  LT_2x1 LT1197 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1343:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1194__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1340:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1692_2486_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2504:150
    ._dfc_wire_2112                          (_LT1197__dfc_wire_2112)
  );
  MUX_3x1 MUX1198 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1344:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_13_2484_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2502:138
    ._dfc_wire_2103_2110                     (_MUX1196__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1342:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1798_2485_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2503:150
    ._dfc_wire_2108                          (_MUX1198__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1199 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1345:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1198__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1344:169
    ._dfc_wire_236 (sink__dfc_wire_2847__dfc_wire_4799)
  );
  dup_1x2 dup1200 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1346:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1178__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1324:135
    ._dfc_wire_68_105 (_dup1200__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1200__dfc_wire_68_113)
  );
  dup_1x2 dup1201 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1347:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR81185__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1331:91
    ._dfc_wire_68_105 (_dup1201__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1201__dfc_wire_68_113)
  );
  ADD_2x1 ADD1202 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1348:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_295_2483_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2501:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1201__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1347:116
    ._dfc_wire_100                          (_ADD1202__dfc_wire_100)
  );
  SHR14_1x1 SHR141203 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1349:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1202__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1348:135
    ._dfc_wire_2103 (_SHR141203__dfc_wire_2103)
  );
  dup_1x3 dup1204 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1350:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141203__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1349:97
    ._dfc_wire_2103_2106 (_dup1204__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1204__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1204__dfc_wire_2103_2113)
  );
  GT_2x1 GT1205 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1351:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1204__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1350:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1826_2482_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2500:150
    ._dfc_wire_2105                          (_GT1205__dfc_wire_2105)
  );
  MUX_3x1 MUX1206 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1352:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1205__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1351:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_1_2480_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2498:138
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1827_2481_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2499:150
    ._dfc_wire_2108                          (_MUX1206__dfc_wire_2108)
  );
  LT_2x1 LT1207 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1353:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1204__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1350:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1792_2479_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2497:150
    ._dfc_wire_2112                          (_LT1207__dfc_wire_2112)
  );
  MUX_3x1 MUX1208 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1354:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_81_2477_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2495:138
    ._dfc_wire_2103_2110                     (_MUX1206__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1352:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1876_2478_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2496:150
    ._dfc_wire_2108                          (_MUX1208__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1209 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1355:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1208__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1354:169
    ._dfc_wire_236 (sink__dfc_wire_2869__dfc_wire_4799)
  );
  dup_1x2 dup1210 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1356:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1179__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1325:114
    ._dfc_wire_68_105 (_dup1210__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1210__dfc_wire_68_113)
  );
  dup_1x2 dup1211 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1357:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR81189__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1335:91
    ._dfc_wire_68_105 (_dup1211__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1211__dfc_wire_68_113)
  );
  ADD_2x1 ADD1212 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1358:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_356_2476_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2494:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1211__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1357:116
    ._dfc_wire_100                          (_ADD1212__dfc_wire_100)
  );
  SHR14_1x1 SHR141213 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1359:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1212__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1358:135
    ._dfc_wire_2103 (_SHR141213__dfc_wire_2103)
  );
  dup_1x3 dup1214 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1360:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141213__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1359:97
    ._dfc_wire_2103_2106 (_dup1214__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1214__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1214__dfc_wire_2103_2113)
  );
  GT_2x1 GT1215 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1361:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1214__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1360:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1825_2475_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2493:150
    ._dfc_wire_2105                          (_GT1215__dfc_wire_2105)
  );
  MUX_3x1 MUX1216 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1362:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1215__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1361:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_44_2473_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2491:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1869_2474_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2492:150
    ._dfc_wire_2108                          (_MUX1216__dfc_wire_2108)
  );
  LT_2x1 LT1217 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1363:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1214__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1360:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1791_2472_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2490:150
    ._dfc_wire_2112                          (_LT1217__dfc_wire_2112)
  );
  MUX_3x1 MUX1218 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1364:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_80_2470_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2488:138
    ._dfc_wire_2103_2110                     (_MUX1216__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1362:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1918_2471_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2489:150
    ._dfc_wire_2108                          (_MUX1218__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1219 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1365:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1218__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1364:169
    ._dfc_wire_236 (sink__dfc_wire_2891__dfc_wire_4799)
  );
  dup_1x2 dup1220 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1366:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1175__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1321:114
    ._dfc_wire_68_105 (_dup1220__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1220__dfc_wire_68_113)
  );
  dup_1x2 dup1221 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1367:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1170__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1316:135
    ._dfc_wire_68_105 (_dup1221__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1221__dfc_wire_68_113)
  );
  ADD_2x1 ADD1222 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1368:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1220__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1366:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_103_2469_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2487:146
    ._dfc_wire_100                          (_ADD1222__dfc_wire_100)
  );
  SHR14_1x1 SHR141223 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1369:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1222__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1368:135
    ._dfc_wire_2103 (_SHR141223__dfc_wire_2103)
  );
  dup_1x3 dup1224 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1370:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141223__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1369:97
    ._dfc_wire_2103_2106 (_dup1224__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1224__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1224__dfc_wire_2103_2113)
  );
  GT_2x1 GT1225 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1371:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1224__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1370:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1636_2468_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2486:150
    ._dfc_wire_2105                          (_GT1225__dfc_wire_2105)
  );
  MUX_3x1 MUX1226 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1372:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1225__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1371:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_85_2466_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2484:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1721_2467_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2485:150
    ._dfc_wire_2108                          (_MUX1226__dfc_wire_2108)
  );
  LT_2x1 LT1227 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1373:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1224__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1370:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1602_2465_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2483:150
    ._dfc_wire_2112                          (_LT1227__dfc_wire_2112)
  );
  MUX_3x1 MUX1228 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1374:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_76_2463_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2481:138
    ._dfc_wire_2103_2110                     (_MUX1226__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1372:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1759_2464_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2482:150
    ._dfc_wire_2108                          (_MUX1228__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1229 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1375:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1228__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1374:169
    ._dfc_wire_236 (sink__dfc_wire_2913__dfc_wire_4799)
  );
  SUB_2x1 SUB1230 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1376:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1220__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1366:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_103_2462_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2480:146
    ._dfc_wire_121    (_SUB1230__dfc_wire_121)
  );
  SHR14_1x1 SHR141231 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1377:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1230__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1376:114
    ._dfc_wire_2103 (_SHR141231__dfc_wire_2103)
  );
  dup_1x3 dup1232 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1378:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141231__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1377:97
    ._dfc_wire_2103_2106 (_dup1232__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1232__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1232__dfc_wire_2103_2113)
  );
  GT_2x1 GT1233 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1379:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1232__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1378:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1722_2461_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2479:150
    ._dfc_wire_2105                          (_GT1233__dfc_wire_2105)
  );
  MUX_3x1 MUX1234 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1380:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1233__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1379:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_39_2459_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2477:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1761_2460_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2478:150
    ._dfc_wire_2108                          (_MUX1234__dfc_wire_2108)
  );
  LT_2x1 LT1235 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1381:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1232__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1378:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1688_2458_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2476:150
    ._dfc_wire_2112                          (_LT1235__dfc_wire_2112)
  );
  MUX_3x1 MUX1236 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1382:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_7_2456_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2474:134
    ._dfc_wire_2103_2110                     (_MUX1234__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1380:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1774_2457_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2475:150
    ._dfc_wire_2108                          (_MUX1236__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1237 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1383:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1236__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1382:169
    ._dfc_wire_236 (sink__dfc_wire_2935__dfc_wire_4799)
  );
  SUB_2x1 SUB1238 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1384:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_356_2455_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2473:146
    ._dfc_wire_118    (_dup1211__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1357:116
    ._dfc_wire_121    (_SUB1238__dfc_wire_121)
  );
  SHR14_1x1 SHR141239 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1385:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1238__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1384:114
    ._dfc_wire_2103 (_SHR141239__dfc_wire_2103)
  );
  dup_1x3 dup1240 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1386:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141239__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1385:97
    ._dfc_wire_2103_2106 (_dup1240__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1240__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1240__dfc_wire_2103_2113)
  );
  GT_2x1 GT1241 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1387:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1240__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1386:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1880_2454_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2472:150
    ._dfc_wire_2105                          (_GT1241__dfc_wire_2105)
  );
  MUX_3x1 MUX1242 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1388:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1241__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1387:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_50_2452_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2470:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1930_2453_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2471:150
    ._dfc_wire_2108                          (_MUX1242__dfc_wire_2108)
  );
  LT_2x1 LT1243 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1389:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1240__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1386:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1846_2451_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2469:150
    ._dfc_wire_2112                          (_LT1243__dfc_wire_2112)
  );
  MUX_3x1 MUX1244 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1390:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_20_2449_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2467:138
    ._dfc_wire_2103_2110                     (_MUX1242__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1388:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1941_2450_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2468:150
    ._dfc_wire_2108                          (_MUX1244__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1245 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1391:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1244__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1390:169
    ._dfc_wire_236 (sink__dfc_wire_2957__dfc_wire_4799)
  );
  SUB_2x1 SUB1246 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1392:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_295_2448_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2466:146
    ._dfc_wire_118    (_dup1201__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1347:116
    ._dfc_wire_121    (_SUB1246__dfc_wire_121)
  );
  SHR14_1x1 SHR141247 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1393:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1246__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1392:114
    ._dfc_wire_2103 (_SHR141247__dfc_wire_2103)
  );
  dup_1x3 dup1248 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1394:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141247__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1393:97
    ._dfc_wire_2103_2106 (_dup1248__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1248__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1248__dfc_wire_2103_2113)
  );
  GT_2x1 GT1249 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1395:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1248__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1394:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1915_2447_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2465:150
    ._dfc_wire_2105                          (_GT1249__dfc_wire_2105)
  );
  MUX_3x1 MUX1250 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1396:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1249__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1395:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_57_2445_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2463:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1972_2446_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2464:150
    ._dfc_wire_2108                          (_MUX1250__dfc_wire_2108)
  );
  LT_2x1 LT1251 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1397:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1248__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1394:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1881_2444_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2462:150
    ._dfc_wire_2112                          (_LT1251__dfc_wire_2112)
  );
  MUX_3x1 MUX1252 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1398:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_75_2442_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2460:138
    ._dfc_wire_2103_2110                     (_MUX1250__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1396:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_2017_2443_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2461:150
    ._dfc_wire_2108                          (_MUX1252__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1253 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1399:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1252__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1398:169
    ._dfc_wire_236 (sink__dfc_wire_2979__dfc_wire_4799)
  );
  SUB_2x1 SUB1254 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1400:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_102_2441_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2459:146
    ._dfc_wire_118    (_dup1191__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1337:116
    ._dfc_wire_121    (_SUB1254__dfc_wire_121)
  );
  SHR14_1x1 SHR141255 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1401:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1254__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1400:114
    ._dfc_wire_2103 (_SHR141255__dfc_wire_2103)
  );
  dup_1x3 dup1256 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1402:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141255__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1401:97
    ._dfc_wire_2103_2106 (_dup1256__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1256__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1256__dfc_wire_2103_2113)
  );
  GT_2x1 GT1257 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1403:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1256__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1402:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1761_2440_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2458:150
    ._dfc_wire_2105                          (_GT1257__dfc_wire_2105)
  );
  MUX_3x1 MUX1258 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1404:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1257__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1403:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_27_2438_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2456:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1788_2439_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2457:150
    ._dfc_wire_2108                          (_MUX1258__dfc_wire_2108)
  );
  LT_2x1 LT1259 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1405:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1256__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1402:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1727_2437_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2455:150
    ._dfc_wire_2112                          (_LT1259__dfc_wire_2112)
  );
  MUX_3x1 MUX1260 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1406:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_13_2435_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2453:138
    ._dfc_wire_2103_2110                     (_MUX1258__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1404:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1775_2436_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2454:150
    ._dfc_wire_2108                          (_MUX1260__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1261 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1407:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1260__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1406:169
    ._dfc_wire_236 (sink__dfc_wire_3001__dfc_wire_4799)
  );
  CAST_1x1_16_32 CAST1262 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1408:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST498__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:644:87
    ._dfc_wire_73 (_CAST1262__dfc_wire_73)
  );
  SHL8_1x1 SHL81263 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1409:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1921 (_CAST1262__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1408:88
    ._dfc_wire_1923 (_SHL81263__dfc_wire_1923)
  );
  CAST_1x1_16_32 CAST1264 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1410:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST698__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:844:87
    ._dfc_wire_73 (_CAST1264__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1265 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1411:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST298__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:444:87
    ._dfc_wire_73 (_CAST1265__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1266 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1412:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST198__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:344:87
    ._dfc_wire_73 (_CAST1266__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1267 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1413:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST798__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:944:87
    ._dfc_wire_73 (_CAST1267__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1268 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1414:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST598__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:744:87
    ._dfc_wire_73 (_CAST1268__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1269 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1415:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST398__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:544:87
    ._dfc_wire_73 (_CAST1269__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1270 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1416:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST98__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:244:83
    ._dfc_wire_73 (_CAST1270__dfc_wire_73)
  );
  SHL8_1x1 SHL81271 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1417:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1921 (_CAST1270__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1416:88
    ._dfc_wire_1923 (_SHL81271__dfc_wire_1923)
  );
  ADD_2x1 ADD1272 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1418:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_SHL81271__dfc_wire_1923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1417:93
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_835_2434_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2452:146
    ._dfc_wire_100                          (_ADD1272__dfc_wire_100)
  );
  dup_1x2 dup1273 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1419:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1266__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1412:88
    ._dfc_wire_68_105 (_dup1273__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1273__dfc_wire_68_113)
  );
  dup_1x2 dup1274 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1420:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1267__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1413:88
    ._dfc_wire_68_105 (_dup1274__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1274__dfc_wire_68_113)
  );
  ADD_2x1 ADD1275 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1421:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_3_2433_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2451:138
    .const_fix_32_0_1__0000000000000080_102 (_dup1274__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1420:116
    ._dfc_wire_100                          (_ADD1275__dfc_wire_100)
  );
  MUL_2x1 MUL1276 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1422:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_744_2432_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2450:146
    ._dfc_wire_104                          (_ADD1275__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1421:135
    ._dfc_wire_107                          (_MUL1276__dfc_wire_107)
  );
  ADD_2x1 ADD1277 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1423:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1276__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1422:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_711_2431_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2449:146
    ._dfc_wire_100                          (_ADD1277__dfc_wire_100)
  );
  MUL_2x1 MUL1278 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1424:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_729_2430_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2448:146
    ._dfc_wire_104                          (_dup1273__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1419:116
    ._dfc_wire_107                          (_MUL1278__dfc_wire_107)
  );
  dup_1x2 dup1279 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1425:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1277__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1423:135
    ._dfc_wire_68_105 (_dup1279__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1279__dfc_wire_68_113)
  );
  ADD_2x1 ADD1280 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1426:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1279__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1425:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_80_2429_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2447:142
    ._dfc_wire_100                          (_ADD1280__dfc_wire_100)
  );
  SHR3_1x1 SHR31281 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1427:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_ADD1280__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1426:135
    ._dfc_wire_1968 (_SHR31281__dfc_wire_1968)
  );
  MUL_2x1 MUL1282 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1428:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_776_2428_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2446:146
    ._dfc_wire_104                          (_dup1274__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1420:116
    ._dfc_wire_107                          (_MUL1282__dfc_wire_107)
  );
  SUB_2x1 SUB1283 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1429:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1279__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1425:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_36_2427_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2445:142
    ._dfc_wire_121    (_SUB1283__dfc_wire_121)
  );
  SHR3_1x1 SHR31284 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1430:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1283__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1429:114
    ._dfc_wire_1968 (_SHR31284__dfc_wire_1968)
  );
  dup_1x2 dup1285 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1431:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1268__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1414:88
    ._dfc_wire_68_105 (_dup1285__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1285__dfc_wire_68_113)
  );
  dup_1x2 dup1286 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1432:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1269__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1415:88
    ._dfc_wire_68_105 (_dup1286__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1286__dfc_wire_68_113)
  );
  ADD_2x1 ADD1287 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1433:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1285__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1431:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_9_2426_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2444:138
    ._dfc_wire_100                          (_ADD1287__dfc_wire_100)
  );
  MUL_2x1 MUL1288 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1434:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_781_2425_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2443:146
    ._dfc_wire_104                          (_ADD1287__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1433:135
    ._dfc_wire_107                          (_MUL1288__dfc_wire_107)
  );
  ADD_2x1 ADD1289 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1435:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1288__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1434:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_678_2424_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2442:146
    ._dfc_wire_100                          (_ADD1289__dfc_wire_100)
  );
  MUL_2x1 MUL1290 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1436:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_670_2423_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2441:146
    ._dfc_wire_104                          (_dup1285__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1431:116
    ._dfc_wire_107                          (_MUL1290__dfc_wire_107)
  );
  dup_1x2 dup1291 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1437:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1289__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1435:135
    ._dfc_wire_68_105 (_dup1291__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1291__dfc_wire_68_113)
  );
  SUB_2x1 SUB1292 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1438:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1291__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1437:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_130_2422_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2440:146
    ._dfc_wire_121    (_SUB1292__dfc_wire_121)
  );
  SHR3_1x1 SHR31293 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1439:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1292__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1438:114
    ._dfc_wire_1968 (_SHR31293__dfc_wire_1968)
  );
  MUL_2x1 MUL1294 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1440:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_719_2421_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2439:146
    ._dfc_wire_104                          (_dup1286__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1432:116
    ._dfc_wire_107                          (_MUL1294__dfc_wire_107)
  );
  SUB_2x1 SUB1295 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1441:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1291__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1437:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_71_2420_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2438:142
    ._dfc_wire_121    (_SUB1295__dfc_wire_121)
  );
  SHR3_1x1 SHR31296 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1442:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1295__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1441:114
    ._dfc_wire_1968 (_SHR31296__dfc_wire_1968)
  );
  dup_1x2 dup1297 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1443:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1272__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1418:135
    ._dfc_wire_68_105 (_dup1297__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1297__dfc_wire_68_113)
  );
  dup_1x2 dup1298 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1444:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHL81263__dfc_wire_1923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1409:93
    ._dfc_wire_68_105 (_dup1298__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1298__dfc_wire_68_113)
  );
  ADD_2x1 ADD1299 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1445:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1297__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1443:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_12_2419_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2437:142
    ._dfc_wire_100                          (_ADD1299__dfc_wire_100)
  );
  SUB_2x1 SUB1300 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1446:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1297__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1443:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_12_2418_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2436:142
    ._dfc_wire_121    (_SUB1300__dfc_wire_121)
  );
  dup_1x2 dup1301 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1447:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1265__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1411:88
    ._dfc_wire_68_105 (_dup1301__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1301__dfc_wire_68_113)
  );
  dup_1x2 dup1302 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1448:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1264__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1410:88
    ._dfc_wire_68_105 (_dup1302__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1302__dfc_wire_68_113)
  );
  ADD_2x1 ADD1303 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1449:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1301__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1447:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_161_2417_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2435:146
    ._dfc_wire_100                          (_ADD1303__dfc_wire_100)
  );
  MUL_2x1 MUL1304 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1450:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_869_2416_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2434:146
    ._dfc_wire_104                          (_ADD1303__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1449:135
    ._dfc_wire_107                          (_MUL1304__dfc_wire_107)
  );
  ADD_2x1 ADD1305 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1451:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1304__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1450:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_768_2415_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2433:146
    ._dfc_wire_100                          (_ADD1305__dfc_wire_100)
  );
  MUL_2x1 MUL1306 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1452:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_622_2414_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2432:146
    ._dfc_wire_104                          (_dup1302__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1448:116
    ._dfc_wire_107                          (_MUL1306__dfc_wire_107)
  );
  dup_1x2 dup1307 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1453:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1305__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1451:135
    ._dfc_wire_68_105 (_dup1307__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1307__dfc_wire_68_113)
  );
  SUB_2x1 SUB1308 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1454:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1307__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1453:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_341_2413_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2431:146
    ._dfc_wire_121    (_SUB1308__dfc_wire_121)
  );
  SHR3_1x1 SHR31309 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1455:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1308__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1454:114
    ._dfc_wire_1968 (_SHR31309__dfc_wire_1968)
  );
  MUL_2x1 MUL1310 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1456:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_839_2412_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2430:146
    ._dfc_wire_104                          (_dup1301__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1447:116
    ._dfc_wire_107                          (_MUL1310__dfc_wire_107)
  );
  ADD_2x1 ADD1311 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1457:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1307__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1453:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_175_2411_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2429:146
    ._dfc_wire_100                          (_ADD1311__dfc_wire_100)
  );
  SHR3_1x1 SHR31312 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1458:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_ADD1311__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1457:135
    ._dfc_wire_1968 (_SHR31312__dfc_wire_1968)
  );
  dup_1x2 dup1313 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1459:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31281__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1427:93
    ._dfc_wire_68_105 (_dup1313__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1313__dfc_wire_68_113)
  );
  dup_1x2 dup1314 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1460:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31293__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1439:93
    ._dfc_wire_68_105 (_dup1314__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1314__dfc_wire_68_113)
  );
  ADD_2x1 ADD1315 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1461:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_11_2410_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2428:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1314__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1460:116
    ._dfc_wire_100                          (_ADD1315__dfc_wire_100)
  );
  SUB_2x1 SUB1316 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1462:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_11_2409_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2427:142
    ._dfc_wire_118    (_dup1314__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1460:116
    ._dfc_wire_121    (_SUB1316__dfc_wire_121)
  );
  dup_1x2 dup1317 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1463:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31284__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1430:93
    ._dfc_wire_68_105 (_dup1317__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1317__dfc_wire_68_113)
  );
  dup_1x2 dup1318 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1464:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31296__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1442:93
    ._dfc_wire_68_105 (_dup1318__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1318__dfc_wire_68_113)
  );
  ADD_2x1 ADD1319 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1465:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1317__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1463:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_39_2408_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2426:142
    ._dfc_wire_100                          (_ADD1319__dfc_wire_100)
  );
  SUB_2x1 SUB1320 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1466:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1317__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1463:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_39_2407_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2425:142
    ._dfc_wire_121    (_SUB1320__dfc_wire_121)
  );
  dup_1x2 dup1321 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1467:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1299__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1445:135
    ._dfc_wire_68_105 (_dup1321__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1321__dfc_wire_68_113)
  );
  dup_1x2 dup1322 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1468:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31312__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1458:93
    ._dfc_wire_68_105 (_dup1322__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1322__dfc_wire_68_113)
  );
  ADD_2x1 ADD1323 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1469:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_169_2406_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2424:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1322__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1468:116
    ._dfc_wire_100                          (_ADD1323__dfc_wire_100)
  );
  SUB_2x1 SUB1324 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1470:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_169_2405_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2423:146
    ._dfc_wire_118    (_dup1322__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1468:116
    ._dfc_wire_121    (_SUB1324__dfc_wire_121)
  );
  dup_1x2 dup1325 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1471:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1300__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1446:114
    ._dfc_wire_68_105 (_dup1325__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1325__dfc_wire_68_113)
  );
  dup_1x2 dup1326 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1472:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31309__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1455:93
    ._dfc_wire_68_105 (_dup1326__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1326__dfc_wire_68_113)
  );
  ADD_2x1 ADD1327 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1473:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_288_2404_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2422:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1326__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1472:116
    ._dfc_wire_100                          (_ADD1327__dfc_wire_100)
  );
  SUB_2x1 SUB1328 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1474:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_288_2403_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2421:146
    ._dfc_wire_118    (_dup1326__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1472:116
    ._dfc_wire_121    (_SUB1328__dfc_wire_121)
  );
  dup_1x2 dup1329 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1475:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1316__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1462:114
    ._dfc_wire_68_105 (_dup1329__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1329__dfc_wire_68_113)
  );
  dup_1x2 dup1330 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1476:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1320__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1466:114
    ._dfc_wire_68_105 (_dup1330__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1330__dfc_wire_68_113)
  );
  ADD_2x1 ADD1331 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1477:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1329__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1475:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_11_2402_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2420:142
    ._dfc_wire_100                          (_ADD1331__dfc_wire_100)
  );
  MUL_2x1 MUL1332 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1478:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1149_2401_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2419:150
    ._dfc_wire_104                          (_ADD1331__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1477:135
    ._dfc_wire_107                          (_MUL1332__dfc_wire_107)
  );
  ADD_2x1 ADD1333 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1479:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1332__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1478:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1291_2400_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2418:150
    ._dfc_wire_100                          (_ADD1333__dfc_wire_100)
  );
  SHR8_1x1 SHR81334 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1480:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD1333__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1479:135
    ._dfc_wire_216 (_SHR81334__dfc_wire_216)
  );
  SUB_2x1 SUB1335 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1481:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1329__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1475:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_11_2399_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2417:142
    ._dfc_wire_121    (_SUB1335__dfc_wire_121)
  );
  MUL_2x1 MUL1336 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1482:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1120_2398_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2416:150
    ._dfc_wire_104                          (_SUB1335__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1481:114
    ._dfc_wire_107                          (_MUL1336__dfc_wire_107)
  );
  ADD_2x1 ADD1337 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1483:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1336__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1482:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1293_2397_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2415:150
    ._dfc_wire_100                          (_ADD1337__dfc_wire_100)
  );
  SHR8_1x1 SHR81338 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1484:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD1337__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1483:135
    ._dfc_wire_216 (_SHR81338__dfc_wire_216)
  );
  dup_1x2 dup1339 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1485:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1323__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1469:135
    ._dfc_wire_68_105 (_dup1339__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1339__dfc_wire_68_113)
  );
  dup_1x2 dup1340 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1486:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1315__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1461:135
    ._dfc_wire_68_105 (_dup1340__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1340__dfc_wire_68_113)
  );
  ADD_2x1 ADD1341 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1487:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1339__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1485:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_48_2396_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2414:142
    ._dfc_wire_100                          (_ADD1341__dfc_wire_100)
  );
  SHR14_1x1 SHR141342 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1488:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1341__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1487:135
    ._dfc_wire_2103 (_SHR141342__dfc_wire_2103)
  );
  dup_1x3 dup1343 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1489:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141342__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1488:97
    ._dfc_wire_2103_2106 (_dup1343__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1343__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1343__dfc_wire_2103_2113)
  );
  GT_2x1 GT1344 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1490:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1343__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1489:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1261_2395_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2413:150
    ._dfc_wire_2105                          (_GT1344__dfc_wire_2105)
  );
  MUX_3x1 MUX1345 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1491:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1344__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1490:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_96_2393_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2411:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1357_2394_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2412:150
    ._dfc_wire_2108                          (_MUX1345__dfc_wire_2108)
  );
  LT_2x1 LT1346 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1492:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1343__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1489:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1227_2392_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2410:150
    ._dfc_wire_2112                          (_LT1346__dfc_wire_2112)
  );
  MUX_3x1 MUX1347 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1493:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_101_2390_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2408:142
    ._dfc_wire_2103_2110                     (_MUX1345__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1491:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1410_2391_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2409:150
    ._dfc_wire_2108                          (_MUX1347__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1348 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1494:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1347__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1493:169
    ._dfc_wire_236 (sink__dfc_wire_3211__dfc_wire_4799)
  );
  dup_1x2 dup1349 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1495:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1327__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1473:135
    ._dfc_wire_68_105 (_dup1349__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1349__dfc_wire_68_113)
  );
  dup_1x2 dup1350 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1496:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR81334__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1480:91
    ._dfc_wire_68_105 (_dup1350__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1350__dfc_wire_68_113)
  );
  ADD_2x1 ADD1351 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1497:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_59_2389_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2407:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1350__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1496:116
    ._dfc_wire_100                          (_ADD1351__dfc_wire_100)
  );
  SHR14_1x1 SHR141352 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1498:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1351__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1497:135
    ._dfc_wire_2103 (_SHR141352__dfc_wire_2103)
  );
  dup_1x3 dup1353 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1499:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141352__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1498:97
    ._dfc_wire_2103_2106 (_dup1353__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1353__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1353__dfc_wire_2103_2113)
  );
  GT_2x1 GT1354 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1500:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1353__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1499:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1496_2388_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2406:150
    ._dfc_wire_2105                          (_GT1354__dfc_wire_2105)
  );
  MUX_3x1 MUX1355 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1501:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1354__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1500:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_55_2386_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2404:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1551_2387_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2405:150
    ._dfc_wire_2108                          (_MUX1355__dfc_wire_2108)
  );
  LT_2x1 LT1356 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1502:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1353__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1499:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1462_2385_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2403:150
    ._dfc_wire_2112                          (_LT1356__dfc_wire_2112)
  );
  MUX_3x1 MUX1357 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1503:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_101_2383_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2401:142
    ._dfc_wire_2103_2110                     (_MUX1355__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1501:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1602_2384_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2402:150
    ._dfc_wire_2108                          (_MUX1357__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1358 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1504:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1357__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1503:169
    ._dfc_wire_236 (sink__dfc_wire_3233__dfc_wire_4799)
  );
  dup_1x2 dup1359 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1505:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1328__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1474:114
    ._dfc_wire_68_105 (_dup1359__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1359__dfc_wire_68_113)
  );
  dup_1x2 dup1360 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1506:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR81338__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1484:91
    ._dfc_wire_68_105 (_dup1360__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1360__dfc_wire_68_113)
  );
  ADD_2x1 ADD1361 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1507:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_18_2382_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2400:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1360__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1506:116
    ._dfc_wire_100                          (_ADD1361__dfc_wire_100)
  );
  SHR14_1x1 SHR141362 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1508:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1361__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1507:135
    ._dfc_wire_2103 (_SHR141362__dfc_wire_2103)
  );
  dup_1x3 dup1363 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1509:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141362__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1508:97
    ._dfc_wire_2103_2106 (_dup1363__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1363__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1363__dfc_wire_2103_2113)
  );
  GT_2x1 GT1364 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1510:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1363__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1509:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1463_2381_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2399:150
    ._dfc_wire_2105                          (_GT1364__dfc_wire_2105)
  );
  MUX_3x1 MUX1365 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1511:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1364__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1510:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_56_2379_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2397:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1519_2380_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2398:150
    ._dfc_wire_2108                          (_MUX1365__dfc_wire_2108)
  );
  LT_2x1 LT1366 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1512:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1363__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1509:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1429_2378_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2396:150
    ._dfc_wire_2112                          (_LT1366__dfc_wire_2112)
  );
  MUX_3x1 MUX1367 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1513:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_64_2376_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2394:138
    ._dfc_wire_2103_2110                     (_MUX1365__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1511:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1540_2377_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2395:150
    ._dfc_wire_2108                          (_MUX1367__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1368 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1514:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1367__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1513:169
    ._dfc_wire_236 (sink__dfc_wire_3255__dfc_wire_4799)
  );
  dup_1x2 dup1369 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1515:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1324__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1470:114
    ._dfc_wire_68_105 (_dup1369__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1369__dfc_wire_68_113)
  );
  dup_1x2 dup1370 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1516:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1319__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1465:135
    ._dfc_wire_68_105 (_dup1370__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1370__dfc_wire_68_113)
  );
  ADD_2x1 ADD1371 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1517:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1369__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1515:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_159_2375_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2393:146
    ._dfc_wire_100                          (_ADD1371__dfc_wire_100)
  );
  SHR14_1x1 SHR141372 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1518:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1371__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1517:135
    ._dfc_wire_2103 (_SHR141372__dfc_wire_2103)
  );
  dup_1x3 dup1373 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1519:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141372__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1518:97
    ._dfc_wire_2103_2106 (_dup1373__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1373__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1373__dfc_wire_2103_2113)
  );
  GT_2x1 GT1374 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1520:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1373__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1519:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1360_2374_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2392:150
    ._dfc_wire_2105                          (_GT1374__dfc_wire_2105)
  );
  MUX_3x1 MUX1375 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1521:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1374__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1520:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_31_2372_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2390:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1391_2373_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2391:150
    ._dfc_wire_2108                          (_MUX1375__dfc_wire_2108)
  );
  LT_2x1 LT1376 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1522:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1373__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1519:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1326_2371_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2389:150
    ._dfc_wire_2112                          (_LT1376__dfc_wire_2112)
  );
  MUX_3x1 MUX1377 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1523:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_114_2369_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2387:142
    ._dfc_wire_2103_2110                     (_MUX1375__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1521:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1450_2370_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2388:150
    ._dfc_wire_2108                          (_MUX1377__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1378 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1524:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1377__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1523:169
    ._dfc_wire_236 (sink__dfc_wire_3277__dfc_wire_4799)
  );
  SUB_2x1 SUB1379 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1525:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1369__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1515:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_159_2368_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2386:146
    ._dfc_wire_121    (_SUB1379__dfc_wire_121)
  );
  SHR14_1x1 SHR141380 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1526:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1379__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1525:114
    ._dfc_wire_2103 (_SHR141380__dfc_wire_2103)
  );
  dup_1x3 dup1381 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1527:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141380__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1526:97
    ._dfc_wire_2103_2106 (_dup1381__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1381__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1381__dfc_wire_2103_2113)
  );
  GT_2x1 GT1382 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1528:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1381__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1527:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1394_2367_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2385:150
    ._dfc_wire_2105                          (_GT1382__dfc_wire_2105)
  );
  MUX_3x1 MUX1383 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1529:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1382__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1528:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_55_2365_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2383:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1449_2366_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2384:150
    ._dfc_wire_2108                          (_MUX1383__dfc_wire_2108)
  );
  LT_2x1 LT1384 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1530:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1381__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1527:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1360_2364_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2382:150
    ._dfc_wire_2112                          (_LT1384__dfc_wire_2112)
  );
  MUX_3x1 MUX1385 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1531:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_71_2362_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2380:138
    ._dfc_wire_2103_2110                     (_MUX1383__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1529:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1487_2363_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2381:150
    ._dfc_wire_2108                          (_MUX1385__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1386 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1532:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1385__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1531:169
    ._dfc_wire_236 (sink__dfc_wire_3299__dfc_wire_4799)
  );
  SUB_2x1 SUB1387 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1533:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_18_2361_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2379:142
    ._dfc_wire_118    (_dup1360__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1506:116
    ._dfc_wire_121    (_SUB1387__dfc_wire_121)
  );
  SHR14_1x1 SHR141388 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1534:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1387__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1533:114
    ._dfc_wire_2103 (_SHR141388__dfc_wire_2103)
  );
  dup_1x3 dup1389 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1535:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141388__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1534:97
    ._dfc_wire_2103_2106 (_dup1389__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1389__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1389__dfc_wire_2103_2113)
  );
  GT_2x1 GT1390 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1536:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1389__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1535:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1520_2360_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2378:150
    ._dfc_wire_2105                          (_GT1390__dfc_wire_2105)
  );
  MUX_3x1 MUX1391 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1537:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1390__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1536:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_35_2358_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2376:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1555_2359_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2377:150
    ._dfc_wire_2108                          (_MUX1391__dfc_wire_2108)
  );
  LT_2x1 LT1392 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1538:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1389__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1535:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1486_2357_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2375:150
    ._dfc_wire_2112                          (_LT1392__dfc_wire_2112)
  );
  MUX_3x1 MUX1393 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1539:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_48_2355_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2373:138
    ._dfc_wire_2103_2110                     (_MUX1391__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1537:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1604_2356_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2374:150
    ._dfc_wire_2108                          (_MUX1393__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1394 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1540:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1393__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1539:169
    ._dfc_wire_236 (sink__dfc_wire_3321__dfc_wire_4799)
  );
  SUB_2x1 SUB1395 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1541:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_59_2354_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2372:142
    ._dfc_wire_118    (_dup1350__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1496:116
    ._dfc_wire_121    (_SUB1395__dfc_wire_121)
  );
  SHR14_1x1 SHR141396 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1542:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1395__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1541:114
    ._dfc_wire_2103 (_SHR141396__dfc_wire_2103)
  );
  dup_1x3 dup1397 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1543:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141396__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1542:97
    ._dfc_wire_2103_2106 (_dup1397__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1397__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1397__dfc_wire_2103_2113)
  );
  GT_2x1 GT1398 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1544:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1397__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1543:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1557_2353_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2371:150
    ._dfc_wire_2105                          (_GT1398__dfc_wire_2105)
  );
  MUX_3x1 MUX1399 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1545:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1398__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1544:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_45_2351_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2369:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1602_2352_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2370:150
    ._dfc_wire_2108                          (_MUX1399__dfc_wire_2108)
  );
  LT_2x1 LT1400 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1546:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1397__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1543:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1523_2350_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2368:150
    ._dfc_wire_2112                          (_LT1400__dfc_wire_2112)
  );
  MUX_3x1 MUX1401 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1547:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_43_2348_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2366:138
    ._dfc_wire_2103_2110                     (_MUX1399__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1545:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1626_2349_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2367:150
    ._dfc_wire_2108                          (_MUX1401__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1402 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1548:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1401__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1547:169
    ._dfc_wire_236 (sink__dfc_wire_3343__dfc_wire_4799)
  );
  SUB_2x1 SUB1403 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1549:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1339__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1485:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_48_2347_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2365:142
    ._dfc_wire_121    (_SUB1403__dfc_wire_121)
  );
  SHR14_1x1 SHR141404 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1550:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1403__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1549:114
    ._dfc_wire_2103 (_SHR141404__dfc_wire_2103)
  );
  dup_1x3 dup1405 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1551:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141404__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1550:97
    ._dfc_wire_2103_2106 (_dup1405__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1405__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1405__dfc_wire_2103_2113)
  );
  GT_2x1 GT1406 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1552:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1405__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1551:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1268_2346_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2364:150
    ._dfc_wire_2105                          (_GT1406__dfc_wire_2105)
  );
  MUX_3x1 MUX1407 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1553:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1406__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1552:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_52_2344_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2362:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1320_2345_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2363:150
    ._dfc_wire_2108                          (_MUX1407__dfc_wire_2108)
  );
  LT_2x1 LT1408 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1554:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1405__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1551:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1234_2343_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2361:150
    ._dfc_wire_2112                          (_LT1408__dfc_wire_2112)
  );
  MUX_3x1 MUX1409 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1555:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_55_2341_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2359:138
    ._dfc_wire_2103_2110                     (_MUX1407__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1553:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1306_2342_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2360:150
    ._dfc_wire_2108                          (_MUX1409__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1410 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1556:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1409__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1555:169
    ._dfc_wire_236 (sink__dfc_wire_3365__dfc_wire_4799)
  );
  CAST_1x1_16_32 CAST1411 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1557:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST501__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:647:87
    ._dfc_wire_73 (_CAST1411__dfc_wire_73)
  );
  SHL8_1x1 SHL81412 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1558:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1921 (_CAST1411__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1557:88
    ._dfc_wire_1923 (_SHL81412__dfc_wire_1923)
  );
  CAST_1x1_16_32 CAST1413 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1559:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST701__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:847:87
    ._dfc_wire_73 (_CAST1413__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1414 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1560:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST301__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:447:87
    ._dfc_wire_73 (_CAST1414__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1415 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1561:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST201__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:347:87
    ._dfc_wire_73 (_CAST1415__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1416 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1562:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST801__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:947:87
    ._dfc_wire_73 (_CAST1416__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1417 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1563:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST601__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:747:87
    ._dfc_wire_73 (_CAST1417__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1418 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1564:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST401__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:547:87
    ._dfc_wire_73 (_CAST1418__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1419 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1565:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST101__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:247:87
    ._dfc_wire_73 (_CAST1419__dfc_wire_73)
  );
  SHL8_1x1 SHL81420 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1566:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1921 (_CAST1419__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1565:88
    ._dfc_wire_1923 (_SHL81420__dfc_wire_1923)
  );
  ADD_2x1 ADD1421 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1567:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_SHL81420__dfc_wire_1923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1566:93
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_902_2340_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2358:146
    ._dfc_wire_100                          (_ADD1421__dfc_wire_100)
  );
  dup_1x2 dup1422 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1568:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1415__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1561:88
    ._dfc_wire_68_105 (_dup1422__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1422__dfc_wire_68_113)
  );
  dup_1x2 dup1423 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1569:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1416__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1562:88
    ._dfc_wire_68_105 (_dup1423__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1423__dfc_wire_68_113)
  );
  ADD_2x1 ADD1424 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1570:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_13_2339_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2357:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1423__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1569:116
    ._dfc_wire_100                          (_ADD1424__dfc_wire_100)
  );
  MUL_2x1 MUL1425 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1571:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_772_2338_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2356:146
    ._dfc_wire_104                          (_ADD1424__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1570:135
    ._dfc_wire_107                          (_MUL1425__dfc_wire_107)
  );
  ADD_2x1 ADD1426 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1572:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1425__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1571:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_778_2337_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2355:146
    ._dfc_wire_100                          (_ADD1426__dfc_wire_100)
  );
  MUL_2x1 MUL1427 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1573:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_708_2336_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2354:146
    ._dfc_wire_104                          (_dup1422__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1568:116
    ._dfc_wire_107                          (_MUL1427__dfc_wire_107)
  );
  dup_1x2 dup1428 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1574:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1426__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1572:135
    ._dfc_wire_68_105 (_dup1428__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1428__dfc_wire_68_113)
  );
  ADD_2x1 ADD1429 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1575:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1428__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1574:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_152_2335_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2353:146
    ._dfc_wire_100                          (_ADD1429__dfc_wire_100)
  );
  SHR3_1x1 SHR31430 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1576:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_ADD1429__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1575:135
    ._dfc_wire_1968 (_SHR31430__dfc_wire_1968)
  );
  MUL_2x1 MUL1431 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1577:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_765_2334_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2352:146
    ._dfc_wire_104                          (_dup1423__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1569:116
    ._dfc_wire_107                          (_MUL1431__dfc_wire_107)
  );
  SUB_2x1 SUB1432 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1578:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1428__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1574:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_163_2333_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2351:146
    ._dfc_wire_121    (_SUB1432__dfc_wire_121)
  );
  SHR3_1x1 SHR31433 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1579:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1432__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1578:114
    ._dfc_wire_1968 (_SHR31433__dfc_wire_1968)
  );
  dup_1x2 dup1434 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1580:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1417__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1563:88
    ._dfc_wire_68_105 (_dup1434__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1434__dfc_wire_68_113)
  );
  dup_1x2 dup1435 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1581:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1418__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1564:88
    ._dfc_wire_68_105 (_dup1435__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1435__dfc_wire_68_113)
  );
  ADD_2x1 ADD1436 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1582:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1434__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1580:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_45_2332_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2350:142
    ._dfc_wire_100                          (_ADD1436__dfc_wire_100)
  );
  MUL_2x1 MUL1437 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1583:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_779_2331_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2349:146
    ._dfc_wire_104                          (_ADD1436__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1582:135
    ._dfc_wire_107                          (_MUL1437__dfc_wire_107)
  );
  ADD_2x1 ADD1438 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1584:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1437__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1583:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_666_2330_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2348:146
    ._dfc_wire_100                          (_ADD1438__dfc_wire_100)
  );
  MUL_2x1 MUL1439 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1585:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_668_2329_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2347:146
    ._dfc_wire_104                          (_dup1434__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1580:116
    ._dfc_wire_107                          (_MUL1439__dfc_wire_107)
  );
  dup_1x2 dup1440 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1586:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1438__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1584:135
    ._dfc_wire_68_105 (_dup1440__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1440__dfc_wire_68_113)
  );
  SUB_2x1 SUB1441 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1587:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1440__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1586:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_92_2328_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2346:142
    ._dfc_wire_121    (_SUB1441__dfc_wire_121)
  );
  SHR3_1x1 SHR31442 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1588:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1441__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1587:114
    ._dfc_wire_1968 (_SHR31442__dfc_wire_1968)
  );
  MUL_2x1 MUL1443 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1589:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_681_2327_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2345:146
    ._dfc_wire_104                          (_dup1435__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1581:116
    ._dfc_wire_107                          (_MUL1443__dfc_wire_107)
  );
  SUB_2x1 SUB1444 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1590:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1440__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1586:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_171_2326_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2344:146
    ._dfc_wire_121    (_SUB1444__dfc_wire_121)
  );
  SHR3_1x1 SHR31445 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1591:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1444__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1590:114
    ._dfc_wire_1968 (_SHR31445__dfc_wire_1968)
  );
  dup_1x2 dup1446 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1592:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1421__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1567:135
    ._dfc_wire_68_105 (_dup1446__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1446__dfc_wire_68_113)
  );
  dup_1x2 dup1447 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1593:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHL81412__dfc_wire_1923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1558:93
    ._dfc_wire_68_105 (_dup1447__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1447__dfc_wire_68_113)
  );
  ADD_2x1 ADD1448 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1594:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1446__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1592:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_160_2325_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2343:146
    ._dfc_wire_100                          (_ADD1448__dfc_wire_100)
  );
  SUB_2x1 SUB1449 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1595:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1446__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1592:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_160_2324_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2342:146
    ._dfc_wire_121    (_SUB1449__dfc_wire_121)
  );
  dup_1x2 dup1450 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1596:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1414__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1560:88
    ._dfc_wire_68_105 (_dup1450__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1450__dfc_wire_68_113)
  );
  dup_1x2 dup1451 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1597:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1413__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1559:88
    ._dfc_wire_68_105 (_dup1451__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1451__dfc_wire_68_113)
  );
  ADD_2x1 ADD1452 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1598:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1450__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1596:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_153_2323_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2341:146
    ._dfc_wire_100                          (_ADD1452__dfc_wire_100)
  );
  MUL_2x1 MUL1453 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1599:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_825_2322_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2340:146
    ._dfc_wire_104                          (_ADD1452__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1598:135
    ._dfc_wire_107                          (_MUL1453__dfc_wire_107)
  );
  ADD_2x1 ADD1454 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1600:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1453__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1599:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_732_2321_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2339:146
    ._dfc_wire_100                          (_ADD1454__dfc_wire_100)
  );
  MUL_2x1 MUL1455 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1601:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_644_2320_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2338:146
    ._dfc_wire_104                          (_dup1451__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1597:116
    ._dfc_wire_107                          (_MUL1455__dfc_wire_107)
  );
  dup_1x2 dup1456 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1602:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1454__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1600:135
    ._dfc_wire_68_105 (_dup1456__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1456__dfc_wire_68_113)
  );
  SUB_2x1 SUB1457 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1603:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1456__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1602:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_274_2319_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2337:146
    ._dfc_wire_121    (_SUB1457__dfc_wire_121)
  );
  SHR3_1x1 SHR31458 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1604:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1457__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1603:114
    ._dfc_wire_1968 (_SHR31458__dfc_wire_1968)
  );
  MUL_2x1 MUL1459 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1605:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_853_2318_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2336:146
    ._dfc_wire_104                          (_dup1450__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1596:116
    ._dfc_wire_107                          (_MUL1459__dfc_wire_107)
  );
  ADD_2x1 ADD1460 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1606:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1456__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1602:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_109_2317_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2335:146
    ._dfc_wire_100                          (_ADD1460__dfc_wire_100)
  );
  SHR3_1x1 SHR31461 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1607:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_ADD1460__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1606:135
    ._dfc_wire_1968 (_SHR31461__dfc_wire_1968)
  );
  dup_1x2 dup1462 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1608:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31430__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1576:93
    ._dfc_wire_68_105 (_dup1462__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1462__dfc_wire_68_113)
  );
  dup_1x2 dup1463 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1609:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31442__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1588:93
    ._dfc_wire_68_105 (_dup1463__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1463__dfc_wire_68_113)
  );
  ADD_2x1 ADD1464 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1610:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1462__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1608:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_11_2316_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2334:142
    ._dfc_wire_100                          (_ADD1464__dfc_wire_100)
  );
  SUB_2x1 SUB1465 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1611:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1462__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1608:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_11_2315_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2333:142
    ._dfc_wire_121    (_SUB1465__dfc_wire_121)
  );
  dup_1x2 dup1466 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1612:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31433__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1579:93
    ._dfc_wire_68_105 (_dup1466__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1466__dfc_wire_68_113)
  );
  dup_1x2 dup1467 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1613:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31445__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1591:93
    ._dfc_wire_68_105 (_dup1467__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1467__dfc_wire_68_113)
  );
  ADD_2x1 ADD1468 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1614:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_27_2314_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2332:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1467__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1613:116
    ._dfc_wire_100                          (_ADD1468__dfc_wire_100)
  );
  SUB_2x1 SUB1469 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1615:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_27_2313_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2331:142
    ._dfc_wire_118    (_dup1467__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1613:116
    ._dfc_wire_121    (_SUB1469__dfc_wire_121)
  );
  dup_1x2 dup1470 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1616:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1448__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1594:135
    ._dfc_wire_68_105 (_dup1470__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1470__dfc_wire_68_113)
  );
  dup_1x2 dup1471 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1617:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31461__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1607:93
    ._dfc_wire_68_105 (_dup1471__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1471__dfc_wire_68_113)
  );
  ADD_2x1 ADD1472 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1618:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_119_2312_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2330:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1471__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1617:116
    ._dfc_wire_100                          (_ADD1472__dfc_wire_100)
  );
  SUB_2x1 SUB1473 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1619:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_119_2311_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2329:146
    ._dfc_wire_118    (_dup1471__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1617:116
    ._dfc_wire_121    (_SUB1473__dfc_wire_121)
  );
  dup_1x2 dup1474 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1620:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1449__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1595:114
    ._dfc_wire_68_105 (_dup1474__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1474__dfc_wire_68_113)
  );
  dup_1x2 dup1475 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1621:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31458__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1604:93
    ._dfc_wire_68_105 (_dup1475__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1475__dfc_wire_68_113)
  );
  ADD_2x1 ADD1476 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1622:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_49_2310_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2328:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1475__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1621:116
    ._dfc_wire_100                          (_ADD1476__dfc_wire_100)
  );
  SUB_2x1 SUB1477 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1623:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_49_2309_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2327:142
    ._dfc_wire_118    (_dup1475__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1621:116
    ._dfc_wire_121    (_SUB1477__dfc_wire_121)
  );
  dup_1x2 dup1478 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1624:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1465__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1611:114
    ._dfc_wire_68_105 (_dup1478__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1478__dfc_wire_68_113)
  );
  dup_1x2 dup1479 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1625:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1469__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1615:114
    ._dfc_wire_68_105 (_dup1479__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1479__dfc_wire_68_113)
  );
  ADD_2x1 ADD1480 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1626:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_172_2308_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2326:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1479__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1625:116
    ._dfc_wire_100                          (_ADD1480__dfc_wire_100)
  );
  MUL_2x1 MUL1481 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1627:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1316_2307_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2325:150
    ._dfc_wire_104                          (_ADD1480__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1626:135
    ._dfc_wire_107                          (_MUL1481__dfc_wire_107)
  );
  ADD_2x1 ADD1482 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1628:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1481__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1627:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1391_2306_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2324:150
    ._dfc_wire_100                          (_ADD1482__dfc_wire_100)
  );
  SHR8_1x1 SHR81483 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1629:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD1482__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1628:135
    ._dfc_wire_216 (_SHR81483__dfc_wire_216)
  );
  SUB_2x1 SUB1484 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1630:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_172_2305_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2323:146
    ._dfc_wire_118    (_dup1479__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1625:116
    ._dfc_wire_121    (_SUB1484__dfc_wire_121)
  );
  MUL_2x1 MUL1485 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1631:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1323_2304_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2322:150
    ._dfc_wire_104                          (_SUB1484__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1630:114
    ._dfc_wire_107                          (_MUL1485__dfc_wire_107)
  );
  ADD_2x1 ADD1486 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1632:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1485__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1631:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1488_2303_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2321:150
    ._dfc_wire_100                          (_ADD1486__dfc_wire_100)
  );
  SHR8_1x1 SHR81487 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1633:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD1486__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1632:135
    ._dfc_wire_216 (_SHR81487__dfc_wire_216)
  );
  dup_1x2 dup1488 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1634:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1472__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1618:135
    ._dfc_wire_68_105 (_dup1488__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1488__dfc_wire_68_113)
  );
  dup_1x2 dup1489 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1635:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1464__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1610:135
    ._dfc_wire_68_105 (_dup1489__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1489__dfc_wire_68_113)
  );
  ADD_2x1 ADD1490 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1636:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_6_2302_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2320:138
    .const_fix_32_0_1__0000000000000080_102 (_dup1489__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1635:116
    ._dfc_wire_100                          (_ADD1490__dfc_wire_100)
  );
  SHR14_1x1 SHR141491 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1637:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1490__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1636:135
    ._dfc_wire_2103 (_SHR141491__dfc_wire_2103)
  );
  dup_1x3 dup1492 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1638:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141491__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1637:97
    ._dfc_wire_2103_2106 (_dup1492__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1492__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1492__dfc_wire_2103_2113)
  );
  GT_2x1 GT1493 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1639:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1492__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1638:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1301_2301_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2319:150
    ._dfc_wire_2105                          (_GT1493__dfc_wire_2105)
  );
  MUX_3x1 MUX1494 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1640:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1493__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1639:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_53_2299_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2317:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1354_2300_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2318:150
    ._dfc_wire_2108                          (_MUX1494__dfc_wire_2108)
  );
  LT_2x1 LT1495 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1641:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1492__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1638:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1267_2298_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2316:150
    ._dfc_wire_2112                          (_LT1495__dfc_wire_2112)
  );
  MUX_3x1 MUX1496 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1642:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_63_2296_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2314:138
    ._dfc_wire_2103_2110                     (_MUX1494__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1640:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1341_2297_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2315:150
    ._dfc_wire_2108                          (_MUX1496__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1497 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1643:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1496__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1642:169
    ._dfc_wire_236 (sink__dfc_wire_3575__dfc_wire_4799)
  );
  dup_1x2 dup1498 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1644:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1476__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1622:135
    ._dfc_wire_68_105 (_dup1498__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1498__dfc_wire_68_113)
  );
  dup_1x2 dup1499 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1645:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR81483__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1629:91
    ._dfc_wire_68_105 (_dup1499__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1499__dfc_wire_68_113)
  );
  ADD_2x1 ADD1500 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1646:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_248_2295_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2313:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1499__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1645:116
    ._dfc_wire_100                          (_ADD1500__dfc_wire_100)
  );
  SHR14_1x1 SHR141501 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1647:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1500__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1646:135
    ._dfc_wire_2103 (_SHR141501__dfc_wire_2103)
  );
  dup_1x3 dup1502 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1648:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141501__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1647:97
    ._dfc_wire_2103_2106 (_dup1502__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1502__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1502__dfc_wire_2103_2113)
  );
  GT_2x1 GT1503 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1649:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1502__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1648:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1643_2294_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2312:150
    ._dfc_wire_2105                          (_GT1503__dfc_wire_2105)
  );
  MUX_3x1 MUX1504 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1650:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1503__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1649:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_55_3239_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3257:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1698_3240_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3258:150
    ._dfc_wire_2108                          (_MUX1504__dfc_wire_2108)
  );
  LT_2x1 LT1505 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1651:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1502__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1648:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1609_3237_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3255:150
    ._dfc_wire_2112                          (_LT1505__dfc_wire_2112)
  );
  MUX_3x1 MUX1506 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1652:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_92_3234_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3252:138
    ._dfc_wire_2103_2110                     (_MUX1504__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1650:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1715_3235_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3253:150
    ._dfc_wire_2108                          (_MUX1506__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1507 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1653:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1506__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1652:169
    ._dfc_wire_236 (sink__dfc_wire_3597__dfc_wire_4799)
  );
  dup_1x2 dup1508 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1654:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1477__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1623:114
    ._dfc_wire_68_105 (_dup1508__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1508__dfc_wire_68_113)
  );
  dup_1x2 dup1509 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1655:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR81487__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1633:91
    ._dfc_wire_68_105 (_dup1509__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1509__dfc_wire_68_113)
  );
  ADD_2x1 ADD1510 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1656:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_340_3232_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3250:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1509__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1655:116
    ._dfc_wire_100                          (_ADD1510__dfc_wire_100)
  );
  SHR14_1x1 SHR141511 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1657:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1510__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1656:135
    ._dfc_wire_2103 (_SHR141511__dfc_wire_2103)
  );
  dup_1x3 dup1512 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1658:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141511__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1657:97
    ._dfc_wire_2103_2106 (_dup1512__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1512__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1512__dfc_wire_2103_2113)
  );
  GT_2x1 GT1513 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1659:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1512__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1658:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1770_3199_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3217:150
    ._dfc_wire_2105                          (_GT1513__dfc_wire_2105)
  );
  MUX_3x1 MUX1514 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1660:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1513__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1659:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_16_3197_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3215:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1786_3198_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3216:150
    ._dfc_wire_2108                          (_MUX1514__dfc_wire_2108)
  );
  LT_2x1 LT1515 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1661:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1512__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1658:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1736_3196_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3214:150
    ._dfc_wire_2112                          (_LT1515__dfc_wire_2112)
  );
  MUX_3x1 MUX1516 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1662:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_LT1515__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1661:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_19_3193_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3211:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1774_3194_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3212:150
    ._dfc_wire_2108                          (_MUX1516__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1517 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1663:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1516__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1662:169
    ._dfc_wire_236 (sink__dfc_wire_3619__dfc_wire_4799)
  );
  dup_1x2 dup1518 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1664:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1473__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1619:114
    ._dfc_wire_68_105 (_dup1518__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1518__dfc_wire_68_113)
  );
  dup_1x2 dup1519 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1665:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1468__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1614:135
    ._dfc_wire_68_105 (_dup1519__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1519__dfc_wire_68_113)
  );
  ADD_2x1 ADD1520 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1666:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_23_2293_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2311:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1519__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1665:116
    ._dfc_wire_100                          (_ADD1520__dfc_wire_100)
  );
  SHR14_1x1 SHR141521 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1667:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1520__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1666:135
    ._dfc_wire_2103 (_SHR141521__dfc_wire_2103)
  );
  dup_1x3 dup1522 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1668:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141521__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1667:97
    ._dfc_wire_2103_2106 (_dup1522__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1522__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1522__dfc_wire_2103_2113)
  );
  GT_2x1 GT1523 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1669:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1522__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1668:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1402_2292_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2310:150
    ._dfc_wire_2105                          (_GT1523__dfc_wire_2105)
  );
  MUX_3x1 MUX1524 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1670:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1523__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1669:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_6_2290_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2308:138
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1408_2291_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2309:150
    ._dfc_wire_2108                          (_MUX1524__dfc_wire_2108)
  );
  LT_2x1 LT1525 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1671:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1522__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1668:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1368_2289_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2307:150
    ._dfc_wire_2112                          (_LT1525__dfc_wire_2112)
  );
  MUX_3x1 MUX1526 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1672:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_LT1525__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1671:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_26_2287_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2305:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1449_2288_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2306:150
    ._dfc_wire_2108                          (_MUX1526__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1527 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1673:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1526__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1672:169
    ._dfc_wire_236 (sink__dfc_wire_3641__dfc_wire_4799)
  );
  SUB_2x1 SUB1528 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1674:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_23_3225_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3243:142
    ._dfc_wire_118    (_dup1519__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1665:116
    ._dfc_wire_121    (_SUB1528__dfc_wire_121)
  );
  SHR14_1x1 SHR141529 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1675:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1528__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1674:114
    ._dfc_wire_2103 (_SHR141529__dfc_wire_2103)
  );
  dup_1x3 dup1530 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1676:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141529__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1675:97
    ._dfc_wire_2103_2106 (_dup1530__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1530__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1530__dfc_wire_2103_2113)
  );
  GT_2x1 GT1531 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1677:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1530__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1676:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1411_3222_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3240:150
    ._dfc_wire_2105                          (_GT1531__dfc_wire_2105)
  );
  MUX_3x1 MUX1532 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1678:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1531__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1677:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_6_3220_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3238:138
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1417_3221_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3239:150
    ._dfc_wire_2108                          (_MUX1532__dfc_wire_2108)
  );
  LT_2x1 LT1533 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1679:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1530__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1676:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1377_3218_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3236:150
    ._dfc_wire_2112                          (_LT1533__dfc_wire_2112)
  );
  MUX_3x1 MUX1534 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1680:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_15_3215_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3233:138
    ._dfc_wire_2103_2110                     (_MUX1532__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1678:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1439_3216_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3234:150
    ._dfc_wire_2108                          (_MUX1534__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1535 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1681:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1534__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1680:169
    ._dfc_wire_236 (sink__dfc_wire_3663__dfc_wire_4799)
  );
  SUB_2x1 SUB1536 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1682:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_340_3214_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3232:146
    ._dfc_wire_118    (_dup1509__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1655:116
    ._dfc_wire_121    (_SUB1536__dfc_wire_121)
  );
  SHR14_1x1 SHR141537 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1683:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1536__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1682:114
    ._dfc_wire_2103 (_SHR141537__dfc_wire_2103)
  );
  dup_1x3 dup1538 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1684:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141537__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1683:97
    ._dfc_wire_2103_2106 (_dup1538__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1538__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1538__dfc_wire_2103_2113)
  );
  GT_2x1 GT1539 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1685:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1538__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1684:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1662_2286_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2304:150
    ._dfc_wire_2105                          (_GT1539__dfc_wire_2105)
  );
  MUX_3x1 MUX1540 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1686:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1539__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1685:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_13_2284_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2302:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1675_2285_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2303:150
    ._dfc_wire_2108                          (_MUX1540__dfc_wire_2108)
  );
  LT_2x1 LT1541 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1687:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1538__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1684:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1628_2283_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2301:150
    ._dfc_wire_2112                          (_LT1541__dfc_wire_2112)
  );
  MUX_3x1 MUX1542 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1688:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_25_2281_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2299:138
    ._dfc_wire_2103_2110                     (_MUX1540__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1686:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1691_2282_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2300:150
    ._dfc_wire_2108                          (_MUX1542__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1543 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1689:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1542__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1688:169
    ._dfc_wire_236 (sink__dfc_wire_3685__dfc_wire_4799)
  );
  SUB_2x1 SUB1544 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1690:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_248_2280_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2298:146
    ._dfc_wire_118    (_dup1499__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1645:116
    ._dfc_wire_121    (_SUB1544__dfc_wire_121)
  );
  SHR14_1x1 SHR141545 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1691:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1544__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1690:114
    ._dfc_wire_2103 (_SHR141545__dfc_wire_2103)
  );
  dup_1x3 dup1546 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1692:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141545__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1691:97
    ._dfc_wire_2103_2106 (_dup1546__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1546__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1546__dfc_wire_2103_2113)
  );
  GT_2x1 GT1547 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1693:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1546__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1692:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1666_2279_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2297:150
    ._dfc_wire_2105                          (_GT1547__dfc_wire_2105)
  );
  MUX_3x1 MUX1548 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1694:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1547__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1693:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_75_2277_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2295:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1741_2278_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2296:150
    ._dfc_wire_2108                          (_MUX1548__dfc_wire_2108)
  );
  LT_2x1 LT1549 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1695:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1546__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1692:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1632_2276_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2294:150
    ._dfc_wire_2112                          (_LT1549__dfc_wire_2112)
  );
  MUX_3x1 MUX1550 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1696:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_114_2274_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2292:142
    ._dfc_wire_2103_2110                     (_MUX1548__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1694:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1771_2275_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2293:150
    ._dfc_wire_2108                          (_MUX1550__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1551 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1697:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1550__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1696:169
    ._dfc_wire_236 (sink__dfc_wire_3707__dfc_wire_4799)
  );
  SUB_2x1 SUB1552 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1698:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_6_2273_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2291:138
    ._dfc_wire_118    (_dup1489__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1635:116
    ._dfc_wire_121    (_SUB1552__dfc_wire_121)
  );
  SHR14_1x1 SHR141553 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1699:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1552__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1698:114
    ._dfc_wire_2103 (_SHR141553__dfc_wire_2103)
  );
  dup_1x3 dup1554 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1700:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141553__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1699:97
    ._dfc_wire_2103_2106 (_dup1554__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1554__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1554__dfc_wire_2103_2113)
  );
  GT_2x1 GT1555 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1701:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1554__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1700:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1338_2272_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2290:150
    ._dfc_wire_2105                          (_GT1555__dfc_wire_2105)
  );
  MUX_3x1 MUX1556 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1702:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1555__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1701:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_31_2270_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2288:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1369_2271_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2289:150
    ._dfc_wire_2108                          (_MUX1556__dfc_wire_2108)
  );
  LT_2x1 LT1557 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1703:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1554__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1700:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1304_2269_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2287:150
    ._dfc_wire_2112                          (_LT1557__dfc_wire_2112)
  );
  MUX_3x1 MUX1558 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1704:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_42_2267_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2285:138
    ._dfc_wire_2103_2110                     (_MUX1556__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1702:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1392_2268_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2286:150
    ._dfc_wire_2108                          (_MUX1558__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1559 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1705:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1558__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1704:169
    ._dfc_wire_236 (sink__dfc_wire_3729__dfc_wire_4799)
  );
  CAST_1x1_16_32 CAST1560 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1706:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST504__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:650:87
    ._dfc_wire_73 (_CAST1560__dfc_wire_73)
  );
  SHL8_1x1 SHL81561 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1707:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1921 (_CAST1560__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1706:88
    ._dfc_wire_1923 (_SHL81561__dfc_wire_1923)
  );
  CAST_1x1_16_32 CAST1562 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1708:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST704__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:850:87
    ._dfc_wire_73 (_CAST1562__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1563 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1709:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST304__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:450:87
    ._dfc_wire_73 (_CAST1563__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1564 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1710:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST204__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:350:87
    ._dfc_wire_73 (_CAST1564__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1565 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1711:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST804__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:950:87
    ._dfc_wire_73 (_CAST1565__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1566 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1712:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST604__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:750:87
    ._dfc_wire_73 (_CAST1566__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1567 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1713:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST404__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:550:87
    ._dfc_wire_73 (_CAST1567__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1568 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1714:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST104__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:250:87
    ._dfc_wire_73 (_CAST1568__dfc_wire_73)
  );
  SHL8_1x1 SHL81569 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1715:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1921 (_CAST1568__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1714:88
    ._dfc_wire_1923 (_SHL81569__dfc_wire_1923)
  );
  ADD_2x1 ADD1570 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1716:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_SHL81569__dfc_wire_1923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1715:93
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_923_2266_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2284:146
    ._dfc_wire_100                          (_ADD1570__dfc_wire_100)
  );
  dup_1x2 dup1571 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1717:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1564__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1710:88
    ._dfc_wire_68_105 (_dup1571__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1571__dfc_wire_68_113)
  );
  dup_1x2 dup1572 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1718:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1565__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1711:88
    ._dfc_wire_68_105 (_dup1572__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1572__dfc_wire_68_113)
  );
  ADD_2x1 ADD1573 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1719:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_32_2265_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2283:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1572__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1718:116
    ._dfc_wire_100                          (_ADD1573__dfc_wire_100)
  );
  MUL_2x1 MUL1574 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1720:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_886_2264_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2282:146
    ._dfc_wire_104                          (_ADD1573__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1719:135
    ._dfc_wire_107                          (_MUL1574__dfc_wire_107)
  );
  ADD_2x1 ADD1575 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1721:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1574__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1720:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_838_2263_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2281:146
    ._dfc_wire_100                          (_ADD1575__dfc_wire_100)
  );
  MUL_2x1 MUL1576 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1722:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_837_2262_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2280:146
    ._dfc_wire_104                          (_dup1571__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1717:116
    ._dfc_wire_107                          (_MUL1576__dfc_wire_107)
  );
  dup_1x2 dup1577 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1723:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1575__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1721:135
    ._dfc_wire_68_105 (_dup1577__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1577__dfc_wire_68_113)
  );
  ADD_2x1 ADD1578 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1724:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1577__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1723:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_155_2261_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2279:146
    ._dfc_wire_100                          (_ADD1578__dfc_wire_100)
  );
  SHR3_1x1 SHR31579 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1725:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_ADD1578__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1724:135
    ._dfc_wire_1968 (_SHR31579__dfc_wire_1968)
  );
  MUL_2x1 MUL1580 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1726:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_913_2260_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2278:146
    ._dfc_wire_104                          (_dup1572__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1718:116
    ._dfc_wire_107                          (_MUL1580__dfc_wire_107)
  );
  SUB_2x1 SUB1581 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1727:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1577__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1723:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_130_2259_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2277:146
    ._dfc_wire_121    (_SUB1581__dfc_wire_121)
  );
  SHR3_1x1 SHR31582 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1728:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1581__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1727:114
    ._dfc_wire_1968 (_SHR31582__dfc_wire_1968)
  );
  dup_1x2 dup1583 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1729:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1566__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1712:88
    ._dfc_wire_68_105 (_dup1583__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1583__dfc_wire_68_113)
  );
  dup_1x2 dup1584 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1730:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1567__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1713:88
    ._dfc_wire_68_105 (_dup1584__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1584__dfc_wire_68_113)
  );
  ADD_2x1 ADD1585 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1731:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_29_2258_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2276:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1584__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1730:116
    ._dfc_wire_100                          (_ADD1585__dfc_wire_100)
  );
  MUL_2x1 MUL1586 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1732:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_965_2257_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2275:146
    ._dfc_wire_104                          (_ADD1585__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1731:135
    ._dfc_wire_107                          (_MUL1586__dfc_wire_107)
  );
  ADD_2x1 ADD1587 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1733:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1586__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1732:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_908_2256_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2274:146
    ._dfc_wire_100                          (_ADD1587__dfc_wire_100)
  );
  MUL_2x1 MUL1588 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1734:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_819_2255_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2273:146
    ._dfc_wire_104                          (_dup1583__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1729:116
    ._dfc_wire_107                          (_MUL1588__dfc_wire_107)
  );
  dup_1x2 dup1589 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1735:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1587__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1733:135
    ._dfc_wire_68_105 (_dup1589__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1589__dfc_wire_68_113)
  );
  SUB_2x1 SUB1590 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1736:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1589__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1735:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_67_2254_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2272:142
    ._dfc_wire_121    (_SUB1590__dfc_wire_121)
  );
  SHR3_1x1 SHR31591 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1737:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1590__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1736:114
    ._dfc_wire_1968 (_SHR31591__dfc_wire_1968)
  );
  MUL_2x1 MUL1592 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1738:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_906_2253_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2271:146
    ._dfc_wire_104                          (_dup1584__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1730:116
    ._dfc_wire_107                          (_MUL1592__dfc_wire_107)
  );
  SUB_2x1 SUB1593 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1739:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1589__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1735:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_71_2252_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2270:142
    ._dfc_wire_121    (_SUB1593__dfc_wire_121)
  );
  SHR3_1x1 SHR31594 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1740:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1593__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1739:114
    ._dfc_wire_1968 (_SHR31594__dfc_wire_1968)
  );
  dup_1x2 dup1595 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1741:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1570__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1716:135
    ._dfc_wire_68_105 (_dup1595__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1595__dfc_wire_68_113)
  );
  dup_1x2 dup1596 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1742:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHL81561__dfc_wire_1923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1707:93
    ._dfc_wire_68_105 (_dup1596__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1596__dfc_wire_68_113)
  );
  ADD_2x1 ADD1597 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1743:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1595__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1741:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_7_2251_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2269:138
    ._dfc_wire_100                          (_ADD1597__dfc_wire_100)
  );
  SUB_2x1 SUB1598 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1744:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1595__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1741:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_7_2250_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2268:138
    ._dfc_wire_121    (_SUB1598__dfc_wire_121)
  );
  dup_1x2 dup1599 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1745:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1563__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1709:88
    ._dfc_wire_68_105 (_dup1599__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1599__dfc_wire_68_113)
  );
  dup_1x2 dup1600 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1746:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1562__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1708:88
    ._dfc_wire_68_105 (_dup1600__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1600__dfc_wire_68_113)
  );
  ADD_2x1 ADD1601 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1747:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1599__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1745:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_86_2249_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2267:142
    ._dfc_wire_100                          (_ADD1601__dfc_wire_100)
  );
  MUL_2x1 MUL1602 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1748:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_986_2248_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2266:146
    ._dfc_wire_104                          (_ADD1601__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1747:135
    ._dfc_wire_107                          (_MUL1602__dfc_wire_107)
  );
  ADD_2x1 ADD1603 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1749:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1602__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1748:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_898_2247_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2265:146
    ._dfc_wire_100                          (_ADD1603__dfc_wire_100)
  );
  MUL_2x1 MUL1604 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1750:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_871_2246_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2264:146
    ._dfc_wire_104                          (_dup1600__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1746:116
    ._dfc_wire_107                          (_MUL1604__dfc_wire_107)
  );
  dup_1x2 dup1605 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1751:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1603__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1749:135
    ._dfc_wire_68_105 (_dup1605__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1605__dfc_wire_68_113)
  );
  SUB_2x1 SUB1606 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1752:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1605__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1751:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_114_2245_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2263:146
    ._dfc_wire_121    (_SUB1606__dfc_wire_121)
  );
  SHR3_1x1 SHR31607 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1753:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1606__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1752:114
    ._dfc_wire_1968 (_SHR31607__dfc_wire_1968)
  );
  MUL_2x1 MUL1608 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1754:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1013_2244_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2262:150
    ._dfc_wire_104                          (_dup1599__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1745:116
    ._dfc_wire_107                          (_MUL1608__dfc_wire_107)
  );
  ADD_2x1 ADD1609 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1755:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1605__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1751:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_17_2243_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2261:142
    ._dfc_wire_100                          (_ADD1609__dfc_wire_100)
  );
  SHR3_1x1 SHR31610 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1756:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_ADD1609__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1755:135
    ._dfc_wire_1968 (_SHR31610__dfc_wire_1968)
  );
  dup_1x2 dup1611 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1757:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31579__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1725:93
    ._dfc_wire_68_105 (_dup1611__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1611__dfc_wire_68_113)
  );
  dup_1x2 dup1612 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1758:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31591__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1737:93
    ._dfc_wire_68_105 (_dup1612__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1612__dfc_wire_68_113)
  );
  ADD_2x1 ADD1613 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1759:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1611__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1757:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_145_2242_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2260:146
    ._dfc_wire_100                          (_ADD1613__dfc_wire_100)
  );
  SUB_2x1 SUB1614 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1760:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1611__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1757:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_145_2241_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2259:146
    ._dfc_wire_121    (_SUB1614__dfc_wire_121)
  );
  dup_1x2 dup1615 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1761:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31582__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1728:93
    ._dfc_wire_68_105 (_dup1615__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1615__dfc_wire_68_113)
  );
  dup_1x2 dup1616 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1762:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31594__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1740:93
    ._dfc_wire_68_105 (_dup1616__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1616__dfc_wire_68_113)
  );
  ADD_2x1 ADD1617 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1763:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1615__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1761:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_71_2240_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2258:142
    ._dfc_wire_100                          (_ADD1617__dfc_wire_100)
  );
  SUB_2x1 SUB1618 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1764:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1615__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1761:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_71_2239_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2257:142
    ._dfc_wire_121    (_SUB1618__dfc_wire_121)
  );
  dup_1x2 dup1619 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1765:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1597__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1743:135
    ._dfc_wire_68_105 (_dup1619__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1619__dfc_wire_68_113)
  );
  dup_1x2 dup1620 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1766:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31610__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1756:93
    ._dfc_wire_68_105 (_dup1620__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1620__dfc_wire_68_113)
  );
  ADD_2x1 ADD1621 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1767:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_65_2238_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2256:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1620__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1766:116
    ._dfc_wire_100                          (_ADD1621__dfc_wire_100)
  );
  SUB_2x1 SUB1622 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1768:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_65_2237_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2255:142
    ._dfc_wire_118    (_dup1620__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1766:116
    ._dfc_wire_121    (_SUB1622__dfc_wire_121)
  );
  dup_1x2 dup1623 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1769:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1598__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1744:114
    ._dfc_wire_68_105 (_dup1623__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1623__dfc_wire_68_113)
  );
  dup_1x2 dup1624 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1770:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31607__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1753:93
    ._dfc_wire_68_105 (_dup1624__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1624__dfc_wire_68_113)
  );
  ADD_2x1 ADD1625 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1771:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_102_2236_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2254:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1624__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1770:116
    ._dfc_wire_100                          (_ADD1625__dfc_wire_100)
  );
  SUB_2x1 SUB1626 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1772:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_102_2235_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2253:146
    ._dfc_wire_118    (_dup1624__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1770:116
    ._dfc_wire_121    (_SUB1626__dfc_wire_121)
  );
  dup_1x2 dup1627 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1773:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1614__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1760:114
    ._dfc_wire_68_105 (_dup1627__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1627__dfc_wire_68_113)
  );
  dup_1x2 dup1628 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1774:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1618__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1764:114
    ._dfc_wire_68_105 (_dup1628__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1628__dfc_wire_68_113)
  );
  ADD_2x1 ADD1629 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1775:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_21_2234_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2252:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1628__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1774:116
    ._dfc_wire_100                          (_ADD1629__dfc_wire_100)
  );
  MUL_2x1 MUL1630 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1776:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1365_2233_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2251:150
    ._dfc_wire_104                          (_ADD1629__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1775:135
    ._dfc_wire_107                          (_MUL1630__dfc_wire_107)
  );
  ADD_2x1 ADD1631 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1777:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1630__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1776:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1478_2232_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2250:150
    ._dfc_wire_100                          (_ADD1631__dfc_wire_100)
  );
  SHR8_1x1 SHR81632 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1778:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD1631__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1777:135
    ._dfc_wire_216 (_SHR81632__dfc_wire_216)
  );
  SUB_2x1 SUB1633 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1779:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_21_2231_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2249:142
    ._dfc_wire_118    (_dup1628__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1774:116
    ._dfc_wire_121    (_SUB1633__dfc_wire_121)
  );
  MUL_2x1 MUL1634 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1780:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1421_2230_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2248:150
    ._dfc_wire_104                          (_SUB1633__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1779:114
    ._dfc_wire_107                          (_MUL1634__dfc_wire_107)
  );
  ADD_2x1 ADD1635 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1781:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1634__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1780:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1561_2229_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2247:150
    ._dfc_wire_100                          (_ADD1635__dfc_wire_100)
  );
  SHR8_1x1 SHR81636 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1782:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD1635__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1781:135
    ._dfc_wire_216 (_SHR81636__dfc_wire_216)
  );
  dup_1x2 dup1637 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1783:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1621__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1767:135
    ._dfc_wire_68_105 (_dup1637__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1637__dfc_wire_68_113)
  );
  dup_1x2 dup1638 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1784:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1613__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1759:135
    ._dfc_wire_68_105 (_dup1638__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1638__dfc_wire_68_113)
  );
  ADD_2x1 ADD1639 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1785:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_52_2228_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2246:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1638__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1784:116
    ._dfc_wire_100                          (_ADD1639__dfc_wire_100)
  );
  SHR14_1x1 SHR141640 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1786:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1639__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1785:135
    ._dfc_wire_2103 (_SHR141640__dfc_wire_2103)
  );
  dup_1x3 dup1641 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1787:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141640__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1786:97
    ._dfc_wire_2103_2106 (_dup1641__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1641__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1641__dfc_wire_2103_2113)
  );
  GT_2x1 GT1642 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1788:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1641__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1787:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1517_2227_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2245:150
    ._dfc_wire_2105                          (_GT1642__dfc_wire_2105)
  );
  MUX_3x1 MUX1643 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1789:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1642__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1788:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_62_2225_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2243:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1579_2226_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2244:150
    ._dfc_wire_2108                          (_MUX1643__dfc_wire_2108)
  );
  LT_2x1 LT1644 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1790:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1641__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1787:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1483_2224_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2242:150
    ._dfc_wire_2112                          (_LT1644__dfc_wire_2112)
  );
  MUX_3x1 MUX1645 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1791:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_92_2222_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2240:138
    ._dfc_wire_2103_2110                     (_MUX1643__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1789:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1612_2223_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2241:150
    ._dfc_wire_2108                          (_MUX1645__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1646 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1792:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1645__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1791:169
    ._dfc_wire_236 (sink__dfc_wire_3939__dfc_wire_4799)
  );
  dup_1x2 dup1647 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1793:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1625__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1771:135
    ._dfc_wire_68_105 (_dup1647__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1647__dfc_wire_68_113)
  );
  dup_1x2 dup1648 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1794:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR81632__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1778:91
    ._dfc_wire_68_105 (_dup1648__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1648__dfc_wire_68_113)
  );
  ADD_2x1 ADD1649 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1795:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_373_2221_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2239:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1648__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1794:116
    ._dfc_wire_100                          (_ADD1649__dfc_wire_100)
  );
  SHR14_1x1 SHR141650 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1796:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1649__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1795:135
    ._dfc_wire_2103 (_SHR141650__dfc_wire_2103)
  );
  dup_1x3 dup1651 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1797:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141650__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1796:97
    ._dfc_wire_2103_2106 (_dup1651__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1651__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1651__dfc_wire_2103_2113)
  );
  GT_2x1 GT1652 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1798:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1651__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1797:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1756_2220_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2238:150
    ._dfc_wire_2105                          (_GT1652__dfc_wire_2105)
  );
  MUX_3x1 MUX1653 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1799:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1652__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1798:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_19_2218_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2236:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1775_2219_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2237:150
    ._dfc_wire_2108                          (_MUX1653__dfc_wire_2108)
  );
  LT_2x1 LT1654 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1800:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1651__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1797:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1722_2217_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2235:150
    ._dfc_wire_2112                          (_LT1654__dfc_wire_2112)
  );
  MUX_3x1 MUX1655 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1801:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_5_2215_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2233:134
    ._dfc_wire_2103_2110                     (_MUX1653__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1799:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1790_2216_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2234:150
    ._dfc_wire_2108                          (_MUX1655__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1656 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1802:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1655__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1801:169
    ._dfc_wire_236 (sink__dfc_wire_3961__dfc_wire_4799)
  );
  dup_1x2 dup1657 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1803:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1626__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1772:114
    ._dfc_wire_68_105 (_dup1657__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1657__dfc_wire_68_113)
  );
  dup_1x2 dup1658 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1804:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR81636__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1782:91
    ._dfc_wire_68_105 (_dup1658__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1658__dfc_wire_68_113)
  );
  ADD_2x1 ADD1659 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1805:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_388_2214_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2232:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1658__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1804:116
    ._dfc_wire_100                          (_ADD1659__dfc_wire_100)
  );
  SHR14_1x1 SHR141660 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1806:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1659__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1805:135
    ._dfc_wire_2103 (_SHR141660__dfc_wire_2103)
  );
  dup_1x3 dup1661 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1807:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141660__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1806:97
    ._dfc_wire_2103_2106 (_dup1661__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1661__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1661__dfc_wire_2103_2113)
  );
  GT_2x1 GT1662 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1808:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1661__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1807:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1763_2213_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2231:150
    ._dfc_wire_2105                          (_GT1662__dfc_wire_2105)
  );
  MUX_3x1 MUX1663 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1809:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1662__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1808:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_41_2211_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2229:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1804_2212_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2230:150
    ._dfc_wire_2108                          (_MUX1663__dfc_wire_2108)
  );
  LT_2x1 LT1664 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1810:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1661__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1807:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1729_2210_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2228:150
    ._dfc_wire_2112                          (_LT1664__dfc_wire_2112)
  );
  MUX_3x1 MUX1665 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1811:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_86_2208_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2226:138
    ._dfc_wire_2103_2110                     (_MUX1663__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1809:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1848_2209_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2227:150
    ._dfc_wire_2108                          (_MUX1665__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1666 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1812:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1665__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1811:169
    ._dfc_wire_236 (sink__dfc_wire_3983__dfc_wire_4799)
  );
  dup_1x2 dup1667 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1813:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1622__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1768:114
    ._dfc_wire_68_105 (_dup1667__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1667__dfc_wire_68_113)
  );
  dup_1x2 dup1668 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1814:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1617__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1763:135
    ._dfc_wire_68_105 (_dup1668__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1668__dfc_wire_68_113)
  );
  ADD_2x1 ADD1669 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1815:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_84_2207_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2225:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1668__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1814:116
    ._dfc_wire_100                          (_ADD1669__dfc_wire_100)
  );
  SHR14_1x1 SHR141670 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1816:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1669__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1815:135
    ._dfc_wire_2103 (_SHR141670__dfc_wire_2103)
  );
  dup_1x3 dup1671 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1817:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141670__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1816:97
    ._dfc_wire_2103_2106 (_dup1671__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1671__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1671__dfc_wire_2103_2113)
  );
  GT_2x1 GT1672 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1818:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1671__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1817:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1441_2206_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2224:150
    ._dfc_wire_2105                          (_GT1672__dfc_wire_2105)
  );
  MUX_3x1 MUX1673 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1819:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1672__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1818:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_11_2204_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2222:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1452_2205_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2223:150
    ._dfc_wire_2108                          (_MUX1673__dfc_wire_2108)
  );
  LT_2x1 LT1674 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1820:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1671__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1817:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1407_2203_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2221:150
    ._dfc_wire_2112                          (_LT1674__dfc_wire_2112)
  );
  MUX_3x1 MUX1675 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1821:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_LT1674__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1820:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_26_2201_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2219:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1446_2202_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2220:150
    ._dfc_wire_2108                          (_MUX1675__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1676 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1822:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1675__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1821:169
    ._dfc_wire_236 (sink__dfc_wire_4005__dfc_wire_4799)
  );
  SUB_2x1 SUB1677 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1823:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_84_2200_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2218:142
    ._dfc_wire_118    (_dup1668__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1814:116
    ._dfc_wire_121    (_SUB1677__dfc_wire_121)
  );
  SHR14_1x1 SHR141678 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1824:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1677__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1823:114
    ._dfc_wire_2103 (_SHR141678__dfc_wire_2103)
  );
  dup_1x3 dup1679 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1825:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141678__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1824:97
    ._dfc_wire_2103_2106 (_dup1679__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1679__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1679__dfc_wire_2103_2113)
  );
  GT_2x1 GT1680 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1826:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1679__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1825:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1371_2199_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2217:150
    ._dfc_wire_2105                          (_GT1680__dfc_wire_2105)
  );
  MUX_3x1 MUX1681 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1827:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1680__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1826:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_20_2197_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2215:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1391_2198_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2216:150
    ._dfc_wire_2108                          (_MUX1681__dfc_wire_2108)
  );
  LT_2x1 LT1682 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1828:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1679__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1825:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1337_2196_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2214:150
    ._dfc_wire_2112                          (_LT1682__dfc_wire_2112)
  );
  MUX_3x1 MUX1683 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1829:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_LT1682__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1828:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_29_2194_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2212:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1391_2195_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2213:150
    ._dfc_wire_2108                          (_MUX1683__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1684 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1830:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1683__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1829:169
    ._dfc_wire_236 (sink__dfc_wire_4027__dfc_wire_4799)
  );
  SUB_2x1 SUB1685 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1831:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_388_2193_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2211:146
    ._dfc_wire_118    (_dup1658__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1804:116
    ._dfc_wire_121    (_SUB1685__dfc_wire_121)
  );
  SHR14_1x1 SHR141686 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1832:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1685__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1831:114
    ._dfc_wire_2103 (_SHR141686__dfc_wire_2103)
  );
  dup_1x3 dup1687 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1833:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141686__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1832:97
    ._dfc_wire_2103_2106 (_dup1687__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1687__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1687__dfc_wire_2103_2113)
  );
  GT_2x1 GT1688 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1834:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1687__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1833:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1865_2192_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2210:150
    ._dfc_wire_2105                          (_GT1688__dfc_wire_2105)
  );
  MUX_3x1 MUX1689 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1835:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1688__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1834:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_75_2190_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2208:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1940_2191_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2209:150
    ._dfc_wire_2108                          (_MUX1689__dfc_wire_2108)
  );
  LT_2x1 LT1690 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1836:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1687__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1833:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1831_2189_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2207:150
    ._dfc_wire_2112                          (_LT1690__dfc_wire_2112)
  );
  MUX_3x1 MUX1691 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1837:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_106_2187_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2205:142
    ._dfc_wire_2103_2110                     (_MUX1689__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1835:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1996_2188_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2206:150
    ._dfc_wire_2108                          (_MUX1691__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1692 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1838:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1691__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1837:169
    ._dfc_wire_236 (sink__dfc_wire_4049__dfc_wire_4799)
  );
  SUB_2x1 SUB1693 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1839:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_373_2186_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2204:146
    ._dfc_wire_118    (_dup1648__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1794:116
    ._dfc_wire_121    (_SUB1693__dfc_wire_121)
  );
  SHR14_1x1 SHR141694 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1840:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1693__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1839:114
    ._dfc_wire_2103 (_SHR141694__dfc_wire_2103)
  );
  dup_1x3 dup1695 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1841:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141694__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1840:97
    ._dfc_wire_2103_2106 (_dup1695__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1695__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1695__dfc_wire_2103_2113)
  );
  GT_2x1 GT1696 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1842:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1695__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1841:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1719_2185_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2203:150
    ._dfc_wire_2105                          (_GT1696__dfc_wire_2105)
  );
  MUX_3x1 MUX1697 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1843:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1696__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1842:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_60_2183_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2201:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1779_2184_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2202:150
    ._dfc_wire_2108                          (_MUX1697__dfc_wire_2108)
  );
  LT_2x1 LT1698 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1844:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1695__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1841:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1685_2182_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2200:150
    ._dfc_wire_2112                          (_LT1698__dfc_wire_2112)
  );
  MUX_3x1 MUX1699 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1845:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_60_2180_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2198:138
    ._dfc_wire_2103_2110                     (_MUX1697__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1843:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1812_2181_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2199:150
    ._dfc_wire_2108                          (_MUX1699__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1700 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1846:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1699__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1845:169
    ._dfc_wire_236 (sink__dfc_wire_4071__dfc_wire_4799)
  );
  SUB_2x1 SUB1701 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1847:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_52_2179_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2197:142
    ._dfc_wire_118    (_dup1638__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1784:116
    ._dfc_wire_121    (_SUB1701__dfc_wire_121)
  );
  SHR14_1x1 SHR141702 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1848:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1701__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1847:114
    ._dfc_wire_2103 (_SHR141702__dfc_wire_2103)
  );
  dup_1x3 dup1703 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1849:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141702__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1848:97
    ._dfc_wire_2103_2106 (_dup1703__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1703__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1703__dfc_wire_2103_2113)
  );
  GT_2x1 GT1704 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1850:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1703__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1849:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1535_2178_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2196:150
    ._dfc_wire_2105                          (_GT1704__dfc_wire_2105)
  );
  MUX_3x1 MUX1705 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1851:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1704__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1850:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_13_2176_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2194:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1548_2177_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2195:150
    ._dfc_wire_2108                          (_MUX1705__dfc_wire_2108)
  );
  LT_2x1 LT1706 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1852:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1703__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1849:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1501_2175_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2193:150
    ._dfc_wire_2112                          (_LT1706__dfc_wire_2112)
  );
  MUX_3x1 MUX1707 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1853:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_29_2173_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2191:138
    ._dfc_wire_2103_2110                     (_MUX1705__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1851:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1596_2174_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2192:150
    ._dfc_wire_2108                          (_MUX1707__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1708 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1854:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1707__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1853:169
    ._dfc_wire_236 (sink__dfc_wire_4093__dfc_wire_4799)
  );
  CAST_1x1_16_32 CAST1709 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1855:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST507__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:653:87
    ._dfc_wire_73 (_CAST1709__dfc_wire_73)
  );
  SHL8_1x1 SHL81710 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1856:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1921 (_CAST1709__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1855:88
    ._dfc_wire_1923 (_SHL81710__dfc_wire_1923)
  );
  CAST_1x1_16_32 CAST1711 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1857:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST707__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:853:87
    ._dfc_wire_73 (_CAST1711__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1712 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1858:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST307__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:453:87
    ._dfc_wire_73 (_CAST1712__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1713 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1859:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST207__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:353:87
    ._dfc_wire_73 (_CAST1713__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1714 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1860:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST807__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:953:87
    ._dfc_wire_73 (_CAST1714__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1715 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1861:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST607__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:753:87
    ._dfc_wire_73 (_CAST1715__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1716 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1862:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST407__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:553:87
    ._dfc_wire_73 (_CAST1716__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1717 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1863:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST107__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:253:87
    ._dfc_wire_73 (_CAST1717__dfc_wire_73)
  );
  SHL8_1x1 SHL81718 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1864:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1921 (_CAST1717__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1863:88
    ._dfc_wire_1923 (_SHL81718__dfc_wire_1923)
  );
  ADD_2x1 ADD1719 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1865:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_SHL81718__dfc_wire_1923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1864:93
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_990_2172_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2190:146
    ._dfc_wire_100                          (_ADD1719__dfc_wire_100)
  );
  dup_1x2 dup1720 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1866:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1713__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1859:88
    ._dfc_wire_68_105 (_dup1720__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1720__dfc_wire_68_113)
  );
  dup_1x2 dup1721 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1867:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1714__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1860:88
    ._dfc_wire_68_105 (_dup1721__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1721__dfc_wire_68_113)
  );
  ADD_2x1 ADD1722 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1868:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1720__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1866:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_274_2171_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2189:146
    ._dfc_wire_100                          (_ADD1722__dfc_wire_100)
  );
  MUL_2x1 MUL1723 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1869:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1154_2170_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2188:150
    ._dfc_wire_104                          (_ADD1722__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1868:135
    ._dfc_wire_107                          (_MUL1723__dfc_wire_107)
  );
  ADD_2x1 ADD1724 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1870:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1723__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1869:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1099_2169_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2187:150
    ._dfc_wire_100                          (_ADD1724__dfc_wire_100)
  );
  MUL_2x1 MUL1725 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1871:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1055_2168_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2186:150
    ._dfc_wire_104                          (_dup1720__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1866:116
    ._dfc_wire_107                          (_MUL1725__dfc_wire_107)
  );
  dup_1x2 dup1726 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1872:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1724__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1870:135
    ._dfc_wire_68_105 (_dup1726__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1726__dfc_wire_68_113)
  );
  ADD_2x1 ADD1727 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1873:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1726__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1872:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_194_2167_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2185:146
    ._dfc_wire_100                          (_ADD1727__dfc_wire_100)
  );
  SHR3_1x1 SHR31728 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1874:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_ADD1727__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1873:135
    ._dfc_wire_1968 (_SHR31728__dfc_wire_1968)
  );
  MUL_2x1 MUL1729 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1875:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_825_2166_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2184:146
    ._dfc_wire_104                          (_dup1721__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1867:116
    ._dfc_wire_107                          (_MUL1729__dfc_wire_107)
  );
  SUB_2x1 SUB1730 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1876:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1726__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1872:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_436_2165_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2183:146
    ._dfc_wire_121    (_SUB1730__dfc_wire_121)
  );
  SHR3_1x1 SHR31731 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1877:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1730__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1876:114
    ._dfc_wire_1968 (_SHR31731__dfc_wire_1968)
  );
  dup_1x2 dup1732 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1878:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1715__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1861:88
    ._dfc_wire_68_105 (_dup1732__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1732__dfc_wire_68_113)
  );
  dup_1x2 dup1733 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1879:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1716__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1862:88
    ._dfc_wire_68_105 (_dup1733__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1733__dfc_wire_68_113)
  );
  ADD_2x1 ADD1734 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1880:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_46_2164_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2182:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1733__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1879:116
    ._dfc_wire_100                          (_ADD1734__dfc_wire_100)
  );
  MUL_2x1 MUL1735 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1881:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1041_2163_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2181:150
    ._dfc_wire_104                          (_ADD1734__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1880:135
    ._dfc_wire_107                          (_MUL1735__dfc_wire_107)
  );
  ADD_2x1 ADD1736 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1882:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1735__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1881:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1007_2162_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2180:150
    ._dfc_wire_100                          (_ADD1736__dfc_wire_100)
  );
  MUL_2x1 MUL1737 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1883:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_876_2161_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2179:146
    ._dfc_wire_104                          (_dup1732__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1878:116
    ._dfc_wire_107                          (_MUL1737__dfc_wire_107)
  );
  dup_1x2 dup1738 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1884:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1736__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1882:135
    ._dfc_wire_68_105 (_dup1738__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1738__dfc_wire_68_113)
  );
  SUB_2x1 SUB1739 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1885:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1738__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1884:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_240_2160_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2178:146
    ._dfc_wire_121    (_SUB1739__dfc_wire_121)
  );
  SHR3_1x1 SHR31740 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1886:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1739__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1885:114
    ._dfc_wire_1968 (_SHR31740__dfc_wire_1968)
  );
  MUL_2x1 MUL1741 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1887:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_980_2159_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2177:146
    ._dfc_wire_104                          (_dup1733__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1879:116
    ._dfc_wire_107                          (_MUL1741__dfc_wire_107)
  );
  SUB_2x1 SUB1742 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1888:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1738__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1884:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_147_2158_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2176:146
    ._dfc_wire_121    (_SUB1742__dfc_wire_121)
  );
  SHR3_1x1 SHR31743 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1889:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1742__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1888:114
    ._dfc_wire_1968 (_SHR31743__dfc_wire_1968)
  );
  dup_1x2 dup1744 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1890:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1719__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1865:135
    ._dfc_wire_68_105 (_dup1744__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1744__dfc_wire_68_113)
  );
  dup_1x2 dup1745 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1891:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHL81710__dfc_wire_1923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1856:93
    ._dfc_wire_68_105 (_dup1745__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1745__dfc_wire_68_113)
  );
  ADD_2x1 ADD1746 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1892:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1744__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1890:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_16_2157_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2175:142
    ._dfc_wire_100                          (_ADD1746__dfc_wire_100)
  );
  SUB_2x1 SUB1747 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1893:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1744__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1890:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_16_2156_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2174:142
    ._dfc_wire_121    (_SUB1747__dfc_wire_121)
  );
  dup_1x2 dup1748 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1894:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1712__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1858:88
    ._dfc_wire_68_105 (_dup1748__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1748__dfc_wire_68_113)
  );
  dup_1x2 dup1749 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1895:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1711__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1857:88
    ._dfc_wire_68_105 (_dup1749__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1749__dfc_wire_68_113)
  );
  ADD_2x1 ADD1750 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1896:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1748__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1894:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_156_2155_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2173:146
    ._dfc_wire_100                          (_ADD1750__dfc_wire_100)
  );
  MUL_2x1 MUL1751 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1897:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_962_2154_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2172:146
    ._dfc_wire_104                          (_ADD1750__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1896:135
    ._dfc_wire_107                          (_MUL1751__dfc_wire_107)
  );
  ADD_2x1 ADD1752 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1898:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1751__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1897:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_917_2153_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2171:146
    ._dfc_wire_100                          (_ADD1752__dfc_wire_100)
  );
  MUL_2x1 MUL1753 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1899:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_784_2152_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2170:146
    ._dfc_wire_104                          (_dup1749__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1895:116
    ._dfc_wire_107                          (_MUL1753__dfc_wire_107)
  );
  dup_1x2 dup1754 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1900:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1752__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1898:135
    ._dfc_wire_68_105 (_dup1754__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1754__dfc_wire_68_113)
  );
  SUB_2x1 SUB1755 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1901:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1754__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1900:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_273_2151_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2169:146
    ._dfc_wire_121    (_SUB1755__dfc_wire_121)
  );
  SHR3_1x1 SHR31756 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1902:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1755__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1901:114
    ._dfc_wire_1968 (_SHR31756__dfc_wire_1968)
  );
  MUL_2x1 MUL1757 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1903:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_996_2150_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2168:146
    ._dfc_wire_104                          (_dup1748__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1894:116
    ._dfc_wire_107                          (_MUL1757__dfc_wire_107)
  );
  ADD_2x1 ADD1758 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1904:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1754__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1900:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_130_2851_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2869:146
    ._dfc_wire_100                          (_ADD1758__dfc_wire_100)
  );
  SHR3_1x1 SHR31759 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1905:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_ADD1758__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1904:135
    ._dfc_wire_1968 (_SHR31759__dfc_wire_1968)
  );
  dup_1x2 dup1760 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1906:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31728__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1874:93
    ._dfc_wire_68_105 (_dup1760__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1760__dfc_wire_68_113)
  );
  dup_1x2 dup1761 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1907:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31740__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1886:93
    ._dfc_wire_68_105 (_dup1761__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1761__dfc_wire_68_113)
  );
  ADD_2x1 ADD1762 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1908:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1760__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1906:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_38_2847_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2865:142
    ._dfc_wire_100                          (_ADD1762__dfc_wire_100)
  );
  SUB_2x1 SUB1763 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1909:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1760__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1906:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_38_2845_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2863:142
    ._dfc_wire_121    (_SUB1763__dfc_wire_121)
  );
  dup_1x2 dup1764 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1910:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31731__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1877:93
    ._dfc_wire_68_105 (_dup1764__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1764__dfc_wire_68_113)
  );
  dup_1x2 dup1765 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1911:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31743__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1889:93
    ._dfc_wire_68_105 (_dup1765__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1765__dfc_wire_68_113)
  );
  ADD_2x1 ADD1766 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1912:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_7_2843_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2861:138
    .const_fix_32_0_1__0000000000000080_102 (_dup1765__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1911:116
    ._dfc_wire_100                          (_ADD1766__dfc_wire_100)
  );
  SUB_2x1 SUB1767 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1913:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_7_2841_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2859:138
    ._dfc_wire_118    (_dup1765__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1911:116
    ._dfc_wire_121    (_SUB1767__dfc_wire_121)
  );
  dup_1x2 dup1768 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1914:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1746__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1892:135
    ._dfc_wire_68_105 (_dup1768__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1768__dfc_wire_68_113)
  );
  dup_1x2 dup1769 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1915:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31759__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1905:93
    ._dfc_wire_68_105 (_dup1769__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1769__dfc_wire_68_113)
  );
  ADD_2x1 ADD1770 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1916:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_70_2838_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2856:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1769__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1915:116
    ._dfc_wire_100                          (_ADD1770__dfc_wire_100)
  );
  SUB_2x1 SUB1771 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1917:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_70_2836_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2854:142
    ._dfc_wire_118    (_dup1769__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1915:116
    ._dfc_wire_121    (_SUB1771__dfc_wire_121)
  );
  dup_1x2 dup1772 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1918:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1747__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1893:114
    ._dfc_wire_68_105 (_dup1772__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1772__dfc_wire_68_113)
  );
  dup_1x2 dup1773 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1919:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31756__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1902:93
    ._dfc_wire_68_105 (_dup1773__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1773__dfc_wire_68_113)
  );
  ADD_2x1 ADD1774 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1920:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_76_2833_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2851:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1773__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1919:116
    ._dfc_wire_100                          (_ADD1774__dfc_wire_100)
  );
  SUB_2x1 SUB1775 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1921:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_76_2832_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2850:142
    ._dfc_wire_118    (_dup1773__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1919:116
    ._dfc_wire_121    (_SUB1775__dfc_wire_121)
  );
  dup_1x2 dup1776 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1922:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1763__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1909:114
    ._dfc_wire_68_105 (_dup1776__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1776__dfc_wire_68_113)
  );
  dup_1x2 dup1777 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1923:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1767__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1913:114
    ._dfc_wire_68_105 (_dup1777__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1777__dfc_wire_68_113)
  );
  ADD_2x1 ADD1778 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1924:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1776__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1922:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_59_2829_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2847:142
    ._dfc_wire_100                          (_ADD1778__dfc_wire_100)
  );
  MUL_2x1 MUL1779 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1925:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1500_2828_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2846:150
    ._dfc_wire_104                          (_ADD1778__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1924:135
    ._dfc_wire_107                          (_MUL1779__dfc_wire_107)
  );
  ADD_2x1 ADD1780 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1926:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1779__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1925:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1646_2826_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2844:150
    ._dfc_wire_100                          (_ADD1780__dfc_wire_100)
  );
  SHR8_1x1 SHR81781 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1927:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD1780__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1926:135
    ._dfc_wire_216 (_SHR81781__dfc_wire_216)
  );
  SUB_2x1 SUB1782 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1928:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1776__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1922:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_59_2823_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2841:142
    ._dfc_wire_121    (_SUB1782__dfc_wire_121)
  );
  MUL_2x1 MUL1783 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1929:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1568_2822_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2840:150
    ._dfc_wire_104                          (_SUB1782__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1928:114
    ._dfc_wire_107                          (_MUL1783__dfc_wire_107)
  );
  ADD_2x1 ADD1784 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1930:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1783__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1929:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1685_2820_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2838:150
    ._dfc_wire_100                          (_ADD1784__dfc_wire_100)
  );
  SHR8_1x1 SHR81785 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1931:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD1784__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1930:135
    ._dfc_wire_216 (_SHR81785__dfc_wire_216)
  );
  dup_1x2 dup1786 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1932:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1770__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1916:135
    ._dfc_wire_68_105 (_dup1786__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1786__dfc_wire_68_113)
  );
  dup_1x2 dup1787 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1933:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1762__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1908:135
    ._dfc_wire_68_105 (_dup1787__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1787__dfc_wire_68_113)
  );
  ADD_2x1 ADD1788 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1934:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_158_2817_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2835:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1787__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1933:116
    ._dfc_wire_100                          (_ADD1788__dfc_wire_100)
  );
  SHR14_1x1 SHR141789 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1935:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1788__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1934:135
    ._dfc_wire_2103 (_SHR141789__dfc_wire_2103)
  );
  dup_1x3 dup1790 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1936:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141789__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1935:97
    ._dfc_wire_2103_2106 (_dup1790__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1790__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1790__dfc_wire_2103_2113)
  );
  GT_2x1 GT1791 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1937:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1790__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1936:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1576_2814_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2832:150
    ._dfc_wire_2105                          (_GT1791__dfc_wire_2105)
  );
  MUX_3x1 MUX1792 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1938:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1791__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1937:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_57_2812_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2830:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1633_2813_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2831:150
    ._dfc_wire_2108                          (_MUX1792__dfc_wire_2108)
  );
  LT_2x1 LT1793 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1939:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1790__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1936:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1542_2810_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2828:150
    ._dfc_wire_2112                          (_LT1793__dfc_wire_2112)
  );
  MUX_3x1 MUX1794 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1940:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_53_2807_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2825:138
    ._dfc_wire_2103_2110                     (_MUX1792__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1938:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1657_2808_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2826:150
    ._dfc_wire_2108                          (_MUX1794__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1795 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1941:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1794__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1940:169
    ._dfc_wire_236 (sink__dfc_wire_4303__dfc_wire_4799)
  );
  dup_1x2 dup1796 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1942:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1774__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1920:135
    ._dfc_wire_68_105 (_dup1796__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1796__dfc_wire_68_113)
  );
  dup_1x2 dup1797 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1943:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR81781__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1927:91
    ._dfc_wire_68_105 (_dup1797__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1797__dfc_wire_68_113)
  );
  ADD_2x1 ADD1798 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1944:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_440_2804_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2822:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1797__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1943:116
    ._dfc_wire_100                          (_ADD1798__dfc_wire_100)
  );
  SHR14_1x1 SHR141799 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1945:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1798__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1944:135
    ._dfc_wire_2103 (_SHR141799__dfc_wire_2103)
  );
  dup_1x3 dup1800 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1946:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141799__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1945:97
    ._dfc_wire_2103_2106 (_dup1800__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1800__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1800__dfc_wire_2103_2113)
  );
  GT_2x1 GT1801 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1947:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1800__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1946:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1908_2802_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2820:150
    ._dfc_wire_2105                          (_GT1801__dfc_wire_2105)
  );
  MUX_3x1 MUX1802 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1948:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1801__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1947:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_51_2799_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2817:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1959_2800_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2818:150
    ._dfc_wire_2108                          (_MUX1802__dfc_wire_2108)
  );
  LT_2x1 LT1803 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1949:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1800__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1946:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1874_2798_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2816:150
    ._dfc_wire_2112                          (_LT1803__dfc_wire_2112)
  );
  MUX_3x1 MUX1804 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1950:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_LT1803__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1949:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_19_2796_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2814:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1956_2797_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2815:150
    ._dfc_wire_2108                          (_MUX1804__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1805 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1951:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1804__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1950:169
    ._dfc_wire_236 (sink__dfc_wire_4325__dfc_wire_4799)
  );
  dup_1x2 dup1806 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1952:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1775__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1921:114
    ._dfc_wire_68_105 (_dup1806__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1806__dfc_wire_68_113)
  );
  dup_1x2 dup1807 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1953:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR81785__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1931:91
    ._dfc_wire_68_105 (_dup1807__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1807__dfc_wire_68_113)
  );
  ADD_2x1 ADD1808 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1954:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_445_2792_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2810:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1807__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1953:116
    ._dfc_wire_100                          (_ADD1808__dfc_wire_100)
  );
  SHR14_1x1 SHR141809 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1955:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1808__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1954:135
    ._dfc_wire_2103 (_SHR141809__dfc_wire_2103)
  );
  dup_1x3 dup1810 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1956:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141809__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1955:97
    ._dfc_wire_2103_2106 (_dup1810__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1810__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1810__dfc_wire_2103_2113)
  );
  GT_2x1 GT1811 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1957:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1810__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1956:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1860_2788_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2806:150
    ._dfc_wire_2105                          (_GT1811__dfc_wire_2105)
  );
  MUX_3x1 MUX1812 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1958:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1811__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1957:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_58_2786_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2804:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1918_2787_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2805:150
    ._dfc_wire_2108                          (_MUX1812__dfc_wire_2108)
  );
  LT_2x1 LT1813 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1959:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1810__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1956:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1826_2785_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2803:150
    ._dfc_wire_2112                          (_LT1813__dfc_wire_2112)
  );
  MUX_3x1 MUX1814 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1960:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_18_2783_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2801:138
    ._dfc_wire_2103_2110                     (_MUX1812__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1958:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1912_2784_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2802:150
    ._dfc_wire_2108                          (_MUX1814__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1815 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1961:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1814__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1960:169
    ._dfc_wire_236 (sink__dfc_wire_4347__dfc_wire_4799)
  );
  dup_1x2 dup1816 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1962:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1771__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1917:114
    ._dfc_wire_68_105 (_dup1816__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1816__dfc_wire_68_113)
  );
  dup_1x2 dup1817 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1963:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1766__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1912:135
    ._dfc_wire_68_105 (_dup1817__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1817__dfc_wire_68_113)
  );
  ADD_2x1 ADD1818 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1964:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_207_2781_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2799:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1817__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1963:116
    ._dfc_wire_100                          (_ADD1818__dfc_wire_100)
  );
  SHR14_1x1 SHR141819 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1965:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1818__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1964:135
    ._dfc_wire_2103 (_SHR141819__dfc_wire_2103)
  );
  dup_1x3 dup1820 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1966:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141819__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1965:97
    ._dfc_wire_2103_2106 (_dup1820__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1820__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1820__dfc_wire_2103_2113)
  );
  GT_2x1 GT1821 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1967:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1820__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1966:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1693_2779_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2797:150
    ._dfc_wire_2105                          (_GT1821__dfc_wire_2105)
  );
  MUX_3x1 MUX1822 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1968:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1821__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1967:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_65_2777_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2795:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1758_2778_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2796:150
    ._dfc_wire_2108                          (_MUX1822__dfc_wire_2108)
  );
  LT_2x1 LT1823 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1969:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1820__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1966:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1659_2776_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2794:150
    ._dfc_wire_2112                          (_LT1823__dfc_wire_2112)
  );
  MUX_3x1 MUX1824 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1970:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_79_2774_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2792:138
    ._dfc_wire_2103_2110                     (_MUX1822__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1968:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1808_2775_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2793:150
    ._dfc_wire_2108                          (_MUX1824__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1825 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1971:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1824__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1970:169
    ._dfc_wire_236 (sink__dfc_wire_4369__dfc_wire_4799)
  );
  SUB_2x1 SUB1826 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1972:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_207_2772_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2790:146
    ._dfc_wire_118    (_dup1817__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1963:116
    ._dfc_wire_121    (_SUB1826__dfc_wire_121)
  );
  SHR14_1x1 SHR141827 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1973:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1826__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1972:114
    ._dfc_wire_2103 (_SHR141827__dfc_wire_2103)
  );
  dup_1x3 dup1828 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1974:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141827__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1973:97
    ._dfc_wire_2103_2106 (_dup1828__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1828__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1828__dfc_wire_2103_2113)
  );
  GT_2x1 GT1829 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1975:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1828__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1974:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1727_2771_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2789:150
    ._dfc_wire_2105                          (_GT1829__dfc_wire_2105)
  );
  MUX_3x1 MUX1830 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1976:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1829__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1975:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_54_2768_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2786:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1781_2769_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2787:150
    ._dfc_wire_2108                          (_MUX1830__dfc_wire_2108)
  );
  LT_2x1 LT1831 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1977:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1828__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1974:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1693_2767_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2785:150
    ._dfc_wire_2112                          (_LT1831__dfc_wire_2112)
  );
  MUX_3x1 MUX1832 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1978:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_97_2765_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2783:138
    ._dfc_wire_2103_2110                     (_MUX1830__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1976:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1806_2766_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2784:150
    ._dfc_wire_2108                          (_MUX1832__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1833 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1979:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1832__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1978:169
    ._dfc_wire_236 (sink__dfc_wire_4391__dfc_wire_4799)
  );
  SUB_2x1 SUB1834 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1980:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_445_2763_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2781:146
    ._dfc_wire_118    (_dup1807__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1953:116
    ._dfc_wire_121    (_SUB1834__dfc_wire_121)
  );
  SHR14_1x1 SHR141835 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1981:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1834__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1980:114
    ._dfc_wire_2103 (_SHR141835__dfc_wire_2103)
  );
  dup_1x3 dup1836 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1982:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141835__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1981:97
    ._dfc_wire_2103_2106 (_dup1836__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1836__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1836__dfc_wire_2103_2113)
  );
  GT_2x1 GT1837 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1983:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1836__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1982:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1936_2761_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2779:150
    ._dfc_wire_2105                          (_GT1837__dfc_wire_2105)
  );
  MUX_3x1 MUX1838 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1984:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1837__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1983:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_32_2759_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2777:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1968_2760_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2778:150
    ._dfc_wire_2108                          (_MUX1838__dfc_wire_2108)
  );
  LT_2x1 LT1839 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1985:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1836__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1982:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1902_2757_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2775:150
    ._dfc_wire_2112                          (_LT1839__dfc_wire_2112)
  );
  MUX_3x1 MUX1840 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1986:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_60_2755_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2773:138
    ._dfc_wire_2103_2110                     (_MUX1838__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1984:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1980_2756_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2774:150
    ._dfc_wire_2108                          (_MUX1840__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1841 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1987:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1840__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1986:169
    ._dfc_wire_236 (sink__dfc_wire_4413__dfc_wire_4799)
  );
  SUB_2x1 SUB1842 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1988:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_440_2753_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2771:146
    ._dfc_wire_118    (_dup1797__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1943:116
    ._dfc_wire_121    (_SUB1842__dfc_wire_121)
  );
  SHR14_1x1 SHR141843 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1989:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1842__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1988:114
    ._dfc_wire_2103 (_SHR141843__dfc_wire_2103)
  );
  dup_1x3 dup1844 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1990:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141843__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1989:97
    ._dfc_wire_2103_2106 (_dup1844__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1844__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1844__dfc_wire_2103_2113)
  );
  GT_2x1 GT1845 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1991:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1844__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1990:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1847_2752_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2770:150
    ._dfc_wire_2105                          (_GT1845__dfc_wire_2105)
  );
  MUX_3x1 MUX1846 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1992:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1845__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1991:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_35_2750_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2768:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1882_2751_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2769:150
    ._dfc_wire_2108                          (_MUX1846__dfc_wire_2108)
  );
  LT_2x1 LT1847 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1993:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1844__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1990:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1813_2749_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2767:150
    ._dfc_wire_2112                          (_LT1847__dfc_wire_2112)
  );
  MUX_3x1 MUX1848 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1994:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_8_2747_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2765:134
    ._dfc_wire_2103_2110                     (_MUX1846__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1992:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1899_2748_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2766:150
    ._dfc_wire_2108                          (_MUX1848__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1849 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1995:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1848__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1994:169
    ._dfc_wire_236 (sink__dfc_wire_4435__dfc_wire_4799)
  );
  SUB_2x1 SUB1850 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1996:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_158_2746_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2764:146
    ._dfc_wire_118    (_dup1787__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1933:116
    ._dfc_wire_121    (_SUB1850__dfc_wire_121)
  );
  SHR14_1x1 SHR141851 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1997:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1850__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1996:114
    ._dfc_wire_2103 (_SHR141851__dfc_wire_2103)
  );
  dup_1x3 dup1852 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1998:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141851__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1997:97
    ._dfc_wire_2103_2106 (_dup1852__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1852__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1852__dfc_wire_2103_2113)
  );
  GT_2x1 GT1853 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1999:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1852__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1998:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1583_2745_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2763:150
    ._dfc_wire_2105                          (_GT1853__dfc_wire_2105)
  );
  MUX_3x1 MUX1854 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2000:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1853__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1999:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_41_2743_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2761:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1624_2744_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2762:150
    ._dfc_wire_2108                          (_MUX1854__dfc_wire_2108)
  );
  LT_2x1 LT1855 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2001:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1852__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1998:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1549_2741_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2759:150
    ._dfc_wire_2112                          (_LT1855__dfc_wire_2112)
  );
  MUX_3x1 MUX1856 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2002:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_32_2739_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2757:138
    ._dfc_wire_2103_2110                     (_MUX1854__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2000:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1597_2740_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2758:150
    ._dfc_wire_2108                          (_MUX1856__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1857 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2003:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1856__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2002:169
    ._dfc_wire_236 (sink__dfc_wire_4457__dfc_wire_4799)
  );
  CAST_1x1_16_32 CAST1858 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2004:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST510__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:656:87
    ._dfc_wire_73 (_CAST1858__dfc_wire_73)
  );
  SHL8_1x1 SHL81859 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2005:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1921 (_CAST1858__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2004:88
    ._dfc_wire_1923 (_SHL81859__dfc_wire_1923)
  );
  CAST_1x1_16_32 CAST1860 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2006:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST710__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:856:87
    ._dfc_wire_73 (_CAST1860__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1861 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2007:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST310__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:456:87
    ._dfc_wire_73 (_CAST1861__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1862 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2008:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST210__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:356:87
    ._dfc_wire_73 (_CAST1862__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1863 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2009:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST810__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:956:87
    ._dfc_wire_73 (_CAST1863__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1864 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2010:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST610__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:756:87
    ._dfc_wire_73 (_CAST1864__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1865 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2011:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST410__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:556:87
    ._dfc_wire_73 (_CAST1865__dfc_wire_73)
  );
  CAST_1x1_16_32 CAST1866 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2012:88
    .clock        (clock),
    .reset        (reset),
    ._dfc_wire_4  (_CAST110__dfc_wire_236),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:256:87
    ._dfc_wire_73 (_CAST1866__dfc_wire_73)
  );
  SHL8_1x1 SHL81867 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2013:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1921 (_CAST1866__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2012:88
    ._dfc_wire_1923 (_SHL81867__dfc_wire_1923)
  );
  ADD_2x1 ADD1868 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2014:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_SHL81867__dfc_wire_1923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2013:93
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_765_2730_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2748:146
    ._dfc_wire_100                          (_ADD1868__dfc_wire_100)
  );
  dup_1x2 dup1869 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2015:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1862__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2008:88
    ._dfc_wire_68_105 (_dup1869__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1869__dfc_wire_68_113)
  );
  dup_1x2 dup1870 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2016:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1863__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2009:88
    ._dfc_wire_68_105 (_dup1870__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1870__dfc_wire_68_113)
  );
  ADD_2x1 ADD1871 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2017:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_88_2727_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2745:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1870__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2016:116
    ._dfc_wire_100                          (_ADD1871__dfc_wire_100)
  );
  MUL_2x1 MUL1872 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2018:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_813_2725_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2743:146
    ._dfc_wire_104                          (_ADD1871__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2017:135
    ._dfc_wire_107                          (_MUL1872__dfc_wire_107)
  );
  ADD_2x1 ADD1873 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2019:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1872__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2018:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_805_2723_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2741:146
    ._dfc_wire_100                          (_ADD1873__dfc_wire_100)
  );
  MUL_2x1 MUL1874 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2020:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_647_2722_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2740:146
    ._dfc_wire_104                          (_dup1869__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2015:116
    ._dfc_wire_107                          (_MUL1874__dfc_wire_107)
  );
  dup_1x2 dup1875 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2021:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1873__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2019:135
    ._dfc_wire_68_105 (_dup1875__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1875__dfc_wire_68_113)
  );
  ADD_2x1 ADD1876 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2022:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1875__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2021:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_243_2717_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2735:146
    ._dfc_wire_100                          (_ADD1876__dfc_wire_100)
  );
  SHR3_1x1 SHR31877 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2023:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_ADD1876__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2022:135
    ._dfc_wire_1968 (_SHR31877__dfc_wire_1968)
  );
  MUL_2x1 MUL1878 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2024:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_779_2714_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2732:146
    ._dfc_wire_104                          (_dup1870__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2016:116
    ._dfc_wire_107                          (_MUL1878__dfc_wire_107)
  );
  SUB_2x1 SUB1879 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2025:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1875__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2021:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_119_2711_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2729:146
    ._dfc_wire_121    (_SUB1879__dfc_wire_121)
  );
  SHR3_1x1 SHR31880 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2026:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1879__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2025:114
    ._dfc_wire_1968 (_SHR31880__dfc_wire_1968)
  );
  dup_1x2 dup1881 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2027:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1864__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2010:88
    ._dfc_wire_68_105 (_dup1881__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1881__dfc_wire_68_113)
  );
  dup_1x2 dup1882 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2028:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1865__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2011:88
    ._dfc_wire_68_105 (_dup1882__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1882__dfc_wire_68_113)
  );
  ADD_2x1 ADD1883 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2029:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1881__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2027:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_131_2706_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2724:146
    ._dfc_wire_100                          (_ADD1883__dfc_wire_100)
  );
  MUL_2x1 MUL1884 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2030:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_808_2704_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2722:146
    ._dfc_wire_104                          (_ADD1883__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2029:135
    ._dfc_wire_107                          (_MUL1884__dfc_wire_107)
  );
  ADD_2x1 ADD1885 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2031:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1884__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2030:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_742_2702_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2720:146
    ._dfc_wire_100                          (_ADD1885__dfc_wire_100)
  );
  MUL_2x1 MUL1886 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2032:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_725_2699_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2717:146
    ._dfc_wire_104                          (_dup1881__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2027:116
    ._dfc_wire_107                          (_MUL1886__dfc_wire_107)
  );
  dup_1x2 dup1887 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2033:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1885__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2031:135
    ._dfc_wire_68_105 (_dup1887__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1887__dfc_wire_68_113)
  );
  SUB_2x1 SUB1888 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2034:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1887__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2033:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_176_2695_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2713:146
    ._dfc_wire_121    (_SUB1888__dfc_wire_121)
  );
  SHR3_1x1 SHR31889 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2035:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1888__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2034:114
    ._dfc_wire_1968 (_SHR31889__dfc_wire_1968)
  );
  MUL_2x1 MUL1890 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2036:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_652_2690_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2708:146
    ._dfc_wire_104                          (_dup1882__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2028:116
    ._dfc_wire_107                          (_MUL1890__dfc_wire_107)
  );
  SUB_2x1 SUB1891 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2037:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1887__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2033:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_313_2689_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2707:146
    ._dfc_wire_121    (_SUB1891__dfc_wire_121)
  );
  SHR3_1x1 SHR31892 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2038:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1891__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2037:114
    ._dfc_wire_1968 (_SHR31892__dfc_wire_1968)
  );
  dup_1x2 dup1893 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2039:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1868__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2014:135
    ._dfc_wire_68_105 (_dup1893__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1893__dfc_wire_68_113)
  );
  dup_1x2 dup1894 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2040:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHL81859__dfc_wire_1923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2005:93
    ._dfc_wire_68_105 (_dup1894__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1894__dfc_wire_68_113)
  );
  ADD_2x1 ADD1895 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2041:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_29_2685_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2703:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1894__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2040:116
    ._dfc_wire_100                          (_ADD1895__dfc_wire_100)
  );
  SUB_2x1 SUB1896 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2042:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_29_2683_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2701:142
    ._dfc_wire_118    (_dup1894__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2040:116
    ._dfc_wire_121    (_SUB1896__dfc_wire_121)
  );
  dup_1x2 dup1897 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2043:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1861__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2007:88
    ._dfc_wire_68_105 (_dup1897__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1897__dfc_wire_68_113)
  );
  dup_1x2 dup1898 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2044:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_CAST1860__dfc_wire_73),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2006:88
    ._dfc_wire_68_105 (_dup1898__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1898__dfc_wire_68_113)
  );
  ADD_2x1 ADD1899 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2045:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1897__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2043:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_3_2675_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2693:138
    ._dfc_wire_100                          (_ADD1899__dfc_wire_100)
  );
  MUL_2x1 MUL1900 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2046:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_769_2674_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2692:146
    ._dfc_wire_104                          (_ADD1899__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2045:135
    ._dfc_wire_107                          (_MUL1900__dfc_wire_107)
  );
  ADD_2x1 ADD1901 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2047:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1900__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2046:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_658_2672_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2690:146
    ._dfc_wire_100                          (_ADD1901__dfc_wire_100)
  );
  MUL_2x1 MUL1902 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2048:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_673_2670_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2688:146
    ._dfc_wire_104                          (_dup1898__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2044:116
    ._dfc_wire_107                          (_MUL1902__dfc_wire_107)
  );
  dup_1x2 dup1903 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2049:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1901__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2047:135
    ._dfc_wire_68_105 (_dup1903__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1903__dfc_wire_68_113)
  );
  SUB_2x1 SUB1904 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2050:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1903__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2049:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_195_2668_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2686:146
    ._dfc_wire_121    (_SUB1904__dfc_wire_121)
  );
  SHR3_1x1 SHR31905 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2051:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_SUB1904__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2050:114
    ._dfc_wire_1968 (_SHR31905__dfc_wire_1968)
  );
  MUL_2x1 MUL1906 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2052:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_732_2664_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2682:146
    ._dfc_wire_104                          (_dup1897__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2043:116
    ._dfc_wire_107                          (_MUL1906__dfc_wire_107)
  );
  ADD_2x1 ADD1907 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2053:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1903__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2049:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_174_2660_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2678:146
    ._dfc_wire_100                          (_ADD1907__dfc_wire_100)
  );
  SHR3_1x1 SHR31908 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2054:93
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_1965 (_ADD1907__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2053:135
    ._dfc_wire_1968 (_SHR31908__dfc_wire_1968)
  );
  dup_1x2 dup1909 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2055:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31877__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2023:93
    ._dfc_wire_68_105 (_dup1909__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1909__dfc_wire_68_113)
  );
  dup_1x2 dup1910 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2056:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31889__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2035:93
    ._dfc_wire_68_105 (_dup1910__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1910__dfc_wire_68_113)
  );
  ADD_2x1 ADD1911 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2057:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_3_2652_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2670:138
    .const_fix_32_0_1__0000000000000080_102 (_dup1910__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2056:116
    ._dfc_wire_100                          (_ADD1911__dfc_wire_100)
  );
  SUB_2x1 SUB1912 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2058:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_3_2651_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2669:138
    ._dfc_wire_118    (_dup1910__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2056:116
    ._dfc_wire_121    (_SUB1912__dfc_wire_121)
  );
  dup_1x2 dup1913 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2059:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31880__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2026:93
    ._dfc_wire_68_105 (_dup1913__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1913__dfc_wire_68_113)
  );
  dup_1x2 dup1914 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2060:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31892__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2038:93
    ._dfc_wire_68_105 (_dup1914__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1914__dfc_wire_68_113)
  );
  ADD_2x1 ADD1915 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2061:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_75_2646_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2664:142
    .const_fix_32_0_1__0000000000000080_102 (_dup1914__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2060:116
    ._dfc_wire_100                          (_ADD1915__dfc_wire_100)
  );
  SUB_2x1 SUB1916 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2062:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_75_2645_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2663:142
    ._dfc_wire_118    (_dup1914__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2060:116
    ._dfc_wire_121    (_SUB1916__dfc_wire_121)
  );
  dup_1x2 dup1917 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2063:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1895__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2041:135
    ._dfc_wire_68_105 (_dup1917__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1917__dfc_wire_68_113)
  );
  dup_1x2 dup1918 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2064:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31908__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2054:93
    ._dfc_wire_68_105 (_dup1918__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1918__dfc_wire_68_113)
  );
  ADD_2x1 ADD1919 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2065:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_235_2644_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2662:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1918__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2064:116
    ._dfc_wire_100                          (_ADD1919__dfc_wire_100)
  );
  SUB_2x1 SUB1920 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2066:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_235_2642_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2660:146
    ._dfc_wire_118    (_dup1918__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2064:116
    ._dfc_wire_121    (_SUB1920__dfc_wire_121)
  );
  dup_1x2 dup1921 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2067:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1896__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2042:114
    ._dfc_wire_68_105 (_dup1921__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1921__dfc_wire_68_113)
  );
  dup_1x2 dup1922 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2068:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR31905__dfc_wire_1968),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2051:93
    ._dfc_wire_68_105 (_dup1922__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1922__dfc_wire_68_113)
  );
  ADD_2x1 ADD1923 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2069:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_121_2641_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2659:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1922__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2068:116
    ._dfc_wire_100                          (_ADD1923__dfc_wire_100)
  );
  SUB_2x1 SUB1924 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2070:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_121_2640_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2658:146
    ._dfc_wire_118    (_dup1922__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2068:116
    ._dfc_wire_121    (_SUB1924__dfc_wire_121)
  );
  dup_1x2 dup1925 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2071:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1912__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2058:114
    ._dfc_wire_68_105 (_dup1925__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1925__dfc_wire_68_113)
  );
  dup_1x2 dup1926 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2072:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1916__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2062:114
    ._dfc_wire_68_105 (_dup1926__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1926__dfc_wire_68_113)
  );
  ADD_2x1 ADD1927 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2073:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1925__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2071:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_24_2638_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2656:142
    ._dfc_wire_100                          (_ADD1927__dfc_wire_100)
  );
  MUL_2x1 MUL1928 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2074:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1238_2637_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2655:150
    ._dfc_wire_104                          (_ADD1927__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2073:135
    ._dfc_wire_107                          (_MUL1928__dfc_wire_107)
  );
  ADD_2x1 ADD1929 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2075:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1928__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2074:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1362_2636_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2654:150
    ._dfc_wire_100                          (_ADD1929__dfc_wire_100)
  );
  SHR8_1x1 SHR81930 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2076:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD1929__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2075:135
    ._dfc_wire_216 (_SHR81930__dfc_wire_216)
  );
  SUB_2x1 SUB1931 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2077:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1925__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2071:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_24_2634_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2652:142
    ._dfc_wire_121    (_SUB1931__dfc_wire_121)
  );
  MUL_2x1 MUL1932 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2078:136
    .clock                                  (clock),
    .reset                                  (reset),
    .const_fix_32_0_1__0000000000000235_108 (_delay_fixed_32_0_1_1277_2633_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2651:150
    ._dfc_wire_104                          (_SUB1931__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2077:114
    ._dfc_wire_107                          (_MUL1932__dfc_wire_107)
  );
  ADD_2x1 ADD1933 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2079:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_MUL1932__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2078:136
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_1379_2631_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2649:150
    ._dfc_wire_100                          (_ADD1933__dfc_wire_100)
  );
  SHR8_1x1 SHR81934 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2080:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_213 (_ADD1933__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2079:135
    ._dfc_wire_216 (_SHR81934__dfc_wire_216)
  );
  dup_1x2 dup1935 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2081:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1919__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2065:135
    ._dfc_wire_68_105 (_dup1935__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1935__dfc_wire_68_113)
  );
  dup_1x2 dup1936 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2082:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1911__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2057:135
    ._dfc_wire_68_105 (_dup1936__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1936__dfc_wire_68_113)
  );
  ADD_2x1 ADD1937 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2083:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1935__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2081:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_39_2625_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2643:142
    ._dfc_wire_100                          (_ADD1937__dfc_wire_100)
  );
  SHR14_1x1 SHR141938 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2084:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1937__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2083:135
    ._dfc_wire_2103 (_SHR141938__dfc_wire_2103)
  );
  dup_1x3 dup1939 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2085:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141938__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2084:97
    ._dfc_wire_2103_2106 (_dup1939__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1939__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1939__dfc_wire_2103_2113)
  );
  GT_2x1 GT1940 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2086:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1939__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2085:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1488_2622_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2640:150
    ._dfc_wire_2105                          (_GT1940__dfc_wire_2105)
  );
  MUX_3x1 MUX1941 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2087:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1940__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2086:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_40_2618_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2636:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1528_2619_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2637:150
    ._dfc_wire_2108                          (_MUX1941__dfc_wire_2108)
  );
  LT_2x1 LT1942 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2088:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1939__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2085:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1454_2615_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2633:150
    ._dfc_wire_2112                          (_LT1942__dfc_wire_2112)
  );
  MUX_3x1 MUX1943 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2089:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_52_2611_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2629:138
    ._dfc_wire_2103_2110                     (_MUX1941__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2087:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1575_2612_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2630:150
    ._dfc_wire_2108                          (_MUX1943__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1944 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2090:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1943__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2089:169
    ._dfc_wire_236 (sink__dfc_wire_4667__dfc_wire_4799)
  );
  dup_1x2 dup1945 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2091:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1923__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2069:135
    ._dfc_wire_68_105 (_dup1945__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1945__dfc_wire_68_113)
  );
  dup_1x2 dup1946 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2092:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR81930__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2076:91
    ._dfc_wire_68_105 (_dup1946__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1946__dfc_wire_68_113)
  );
  ADD_2x1 ADD1947 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2093:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_342_2609_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2627:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1946__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2092:116
    ._dfc_wire_100                          (_ADD1947__dfc_wire_100)
  );
  SHR14_1x1 SHR141948 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2094:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1947__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2093:135
    ._dfc_wire_2103 (_SHR141948__dfc_wire_2103)
  );
  dup_1x3 dup1949 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2095:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141948__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2094:97
    ._dfc_wire_2103_2106 (_dup1949__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1949__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1949__dfc_wire_2103_2113)
  );
  GT_2x1 GT1950 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2096:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1949__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2095:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1643_2604_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2622:150
    ._dfc_wire_2105                          (_GT1950__dfc_wire_2105)
  );
  MUX_3x1 MUX1951 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2097:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1950__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2096:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_29_2600_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2618:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1672_2601_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2619:150
    ._dfc_wire_2108                          (_MUX1951__dfc_wire_2108)
  );
  LT_2x1 LT1952 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2098:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1949__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2095:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1609_2599_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2617:150
    ._dfc_wire_2112                          (_LT1952__dfc_wire_2112)
  );
  MUX_3x1 MUX1953 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2099:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_LT1952__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2098:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_62_2596_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2614:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1702_2597_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2615:150
    ._dfc_wire_2108                          (_MUX1953__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1954 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2100:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1953__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2099:169
    ._dfc_wire_236 (sink__dfc_wire_4689__dfc_wire_4799)
  );
  dup_1x2 dup1955 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2101:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1924__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2070:114
    ._dfc_wire_68_105 (_dup1955__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1955__dfc_wire_68_113)
  );
  dup_1x2 dup1956 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2102:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SHR81934__dfc_wire_216),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2080:91
    ._dfc_wire_68_105 (_dup1956__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1956__dfc_wire_68_113)
  );
  ADD_2x1 ADD1957 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2103:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_delay_fixed_32_0_1_346_2591_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2609:146
    .const_fix_32_0_1__0000000000000080_102 (_dup1956__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2102:116
    ._dfc_wire_100                          (_ADD1957__dfc_wire_100)
  );
  SHR14_1x1 SHR141958 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2104:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1957__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2103:135
    ._dfc_wire_2103 (_SHR141958__dfc_wire_2103)
  );
  dup_1x3 dup1959 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2105:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141958__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2104:97
    ._dfc_wire_2103_2106 (_dup1959__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1959__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1959__dfc_wire_2103_2113)
  );
  GT_2x1 GT1960 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2106:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1959__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2105:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1692_2585_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2603:150
    ._dfc_wire_2105                          (_GT1960__dfc_wire_2105)
  );
  MUX_3x1 MUX1961 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2107:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1960__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2106:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_23_2561_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2579:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1715_2562_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2580:150
    ._dfc_wire_2108                          (_MUX1961__dfc_wire_2108)
  );
  LT_2x1 LT1962 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2108:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1959__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2105:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1658_2584_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2602:150
    ._dfc_wire_2112                          (_LT1962__dfc_wire_2112)
  );
  MUX_3x1 MUX1963 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2109:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_LT1962__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2108:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_19_2581_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2599:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1741_2582_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2600:150
    ._dfc_wire_2108                          (_MUX1963__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1964 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2110:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1963__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2109:169
    ._dfc_wire_236 (sink__dfc_wire_4711__dfc_wire_4799)
  );
  dup_1x2 dup1965 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2111:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_SUB1920__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2066:114
    ._dfc_wire_68_105 (_dup1965__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1965__dfc_wire_68_113)
  );
  dup_1x2 dup1966 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2112:116
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_84     (_ADD1915__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2061:135
    ._dfc_wire_68_105 (_dup1966__dfc_wire_68_105),
    ._dfc_wire_68_113 (_dup1966__dfc_wire_68_113)
  );
  ADD_2x1 ADD1967 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2113:135
    .clock                                  (clock),
    .reset                                  (reset),
    ._dfc_wire_98                           (_dup1965__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2111:116
    .const_fix_32_0_1__0000000000000080_102 (_delay_fixed_32_0_1_24_2578_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2596:142
    ._dfc_wire_100                          (_ADD1967__dfc_wire_100)
  );
  SHR14_1x1 SHR141968 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2114:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_ADD1967__dfc_wire_100),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2113:135
    ._dfc_wire_2103 (_SHR141968__dfc_wire_2103)
  );
  dup_1x3 dup1969 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2115:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141968__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2114:97
    ._dfc_wire_2103_2106 (_dup1969__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1969__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1969__dfc_wire_2103_2113)
  );
  GT_2x1 GT1970 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2116:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1969__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2115:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1419_2575_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2593:150
    ._dfc_wire_2105                          (_GT1970__dfc_wire_2105)
  );
  MUX_3x1 MUX1971 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2117:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1970__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2116:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_15_2572_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2590:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1434_2573_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2591:150
    ._dfc_wire_2108                          (_MUX1971__dfc_wire_2108)
  );
  LT_2x1 LT1972 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2118:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1969__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2115:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1385_2571_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2589:150
    ._dfc_wire_2112                          (_LT1972__dfc_wire_2112)
  );
  MUX_3x1 MUX1973 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2119:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_LT1972__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2118:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_6_2568_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2586:138
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1424_2569_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2587:150
    ._dfc_wire_2108                          (_MUX1973__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1974 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2120:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1973__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2119:169
    ._dfc_wire_236 (sink__dfc_wire_4733__dfc_wire_4799)
  );
  SUB_2x1 SUB1975 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2121:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1965__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2111:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_24_2563_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2581:142
    ._dfc_wire_121    (_SUB1975__dfc_wire_121)
  );
  SHR14_1x1 SHR141976 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2122:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1975__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2121:114
    ._dfc_wire_2103 (_SHR141976__dfc_wire_2103)
  );
  dup_1x3 dup1977 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2123:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141976__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2122:97
    ._dfc_wire_2103_2106 (_dup1977__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1977__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1977__dfc_wire_2103_2113)
  );
  GT_2x1 GT1978 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2124:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1977__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2123:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1327_3062_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3080:150
    ._dfc_wire_2105                          (_GT1978__dfc_wire_2105)
  );
  MUX_3x1 MUX1979 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2125:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1978__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2124:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_43_3058_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3076:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1370_3059_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3077:150
    ._dfc_wire_2108                          (_MUX1979__dfc_wire_2108)
  );
  LT_2x1 LT1980 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2126:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1977__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2123:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1293_3056_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3074:150
    ._dfc_wire_2112                          (_LT1980__dfc_wire_2112)
  );
  MUX_3x1 MUX1981 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2127:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_LT1980__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2126:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_26_3052_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3070:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1377_3053_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3071:150
    ._dfc_wire_2108                          (_MUX1981__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1982 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2128:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1981__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2127:169
    ._dfc_wire_236 (sink__dfc_wire_4755__dfc_wire_4799)
  );
  SUB_2x1 SUB1983 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2129:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_346_3048_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3066:146
    ._dfc_wire_118    (_dup1956__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2102:116
    ._dfc_wire_121    (_SUB1983__dfc_wire_121)
  );
  SHR14_1x1 SHR141984 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2130:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1983__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2129:114
    ._dfc_wire_2103 (_SHR141984__dfc_wire_2103)
  );
  dup_1x3 dup1985 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2131:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141984__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2130:97
    ._dfc_wire_2103_2106 (_dup1985__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1985__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1985__dfc_wire_2103_2113)
  );
  GT_2x1 GT1986 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2132:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1985__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2131:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1714_3042_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3060:150
    ._dfc_wire_2105                          (_GT1986__dfc_wire_2105)
  );
  MUX_3x1 MUX1987 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2133:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1986__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2132:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_69_3038_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3056:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1783_3039_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3057:150
    ._dfc_wire_2108                          (_MUX1987__dfc_wire_2108)
  );
  LT_2x1 LT1988 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2134:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1985__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2131:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1680_3035_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3053:150
    ._dfc_wire_2112                          (_LT1988__dfc_wire_2112)
  );
  MUX_3x1 MUX1989 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2135:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_94_3031_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3049:138
    ._dfc_wire_2103_2110                     (_MUX1987__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2133:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1825_3032_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3050:150
    ._dfc_wire_2108                          (_MUX1989__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1990 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2136:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1989__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2135:169
    ._dfc_wire_236 (sink__dfc_wire_4777__dfc_wire_4799)
  );
  SUB_2x1 SUB1991 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2137:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_delay_fixed_32_0_1_342_3228_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3246:146
    ._dfc_wire_118    (_dup1946__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2092:116
    ._dfc_wire_121    (_SUB1991__dfc_wire_121)
  );
  SHR14_1x1 SHR141992 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2138:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1991__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2137:114
    ._dfc_wire_2103 (_SHR141992__dfc_wire_2103)
  );
  dup_1x3 dup1993 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2139:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR141992__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2138:97
    ._dfc_wire_2103_2106 (_dup1993__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup1993__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup1993__dfc_wire_2103_2113)
  );
  GT_2x1 GT1994 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2140:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup1993__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2139:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1711_3024_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3042:150
    ._dfc_wire_2105                          (_GT1994__dfc_wire_2105)
  );
  MUX_3x1 MUX1995 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2141:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT1994__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2140:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_13_3022_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3040:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1724_3023_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3041:150
    ._dfc_wire_2108                          (_MUX1995__dfc_wire_2108)
  );
  LT_2x1 LT1996 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2142:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup1993__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2139:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1677_3020_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3038:150
    ._dfc_wire_2112                          (_LT1996__dfc_wire_2112)
  );
  MUX_3x1 MUX1997 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2143:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_LT1996__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2142:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_9_3016_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3034:138
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1753_3017_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3035:150
    ._dfc_wire_2108                          (_MUX1997__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST1998 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2144:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX1997__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2143:169
    ._dfc_wire_236 (sink__dfc_wire_4799__dfc_wire_4799)
  );
  SUB_2x1 SUB1999 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2145:114
    .clock            (clock),
    .reset            (reset),
    ._dfc_wire_72_122 (_dup1935__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2081:116
    ._dfc_wire_118    (_delay_fixed_32_0_1_39_3013_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3031:142
    ._dfc_wire_121    (_SUB1999__dfc_wire_121)
  );
  SHR14_1x1 SHR142000 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2146:97
    .clock          (clock),
    .reset          (reset),
    ._dfc_wire_2100 (_SUB1999__dfc_wire_121),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2145:114
    ._dfc_wire_2103 (_SHR142000__dfc_wire_2103)
  );
  dup_1x3 dup2001 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2147:154
    .clock               (clock),
    .reset               (reset),
    ._dfc_wire_2103      (_SHR142000__dfc_wire_2103),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2146:97
    ._dfc_wire_2103_2106 (_dup2001__dfc_wire_2103_2106),
    ._dfc_wire_2103_2110 (_dup2001__dfc_wire_2103_2110),
    ._dfc_wire_2103_2113 (_dup2001__dfc_wire_2103_2113)
  );
  GT_2x1 GT2002 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2148:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2106                     (_dup2001__dfc_wire_2103_2106),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2147:154
    .const_fix_32_0_1__00000000000000ff_2107 (_delay_fixed_32_0_1_1455_3008_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3026:150
    ._dfc_wire_2105                          (_GT2002__dfc_wire_2105)
  );
  MUX_3x1 MUX2003 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2149:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_GT2002__dfc_wire_2105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2148:139
    ._dfc_wire_2103_2110                     (_delay_fixed_32_0_1_45_3005_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3023:142
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1500_3006_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3024:150
    ._dfc_wire_2108                          (_MUX2003__dfc_wire_2108)
  );
  LT_2x1 LT2004 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2150:139
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2103_2113                     (_dup2001__dfc_wire_2103_2113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2147:154
    .const_fix_32_0_1__ffffffffffffff00_2114 (_delay_fixed_32_0_1_1421_3003_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3021:150
    ._dfc_wire_2112                          (_LT2004__dfc_wire_2112)
  );
  MUX_3x1 MUX2005 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2151:169
    .clock                                   (clock),
    .reset                                   (reset),
    ._dfc_wire_2105                          (_delay_fixed_1_0_0_25_2999_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3017:138
    ._dfc_wire_2103_2110                     (_MUX2003__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2149:169
    .const_fix_32_0_1__00000000000000ff_2111 (_delay_fixed_32_0_1_1501_3000_out),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3018:150
    ._dfc_wire_2108                          (_MUX2005__dfc_wire_2108)
  );
  CAST_1x1_32_16 CAST2006 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2152:91
    .clock         (clock),
    .reset         (reset),
    ._dfc_wire_234 (_MUX2005__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2151:169
    ._dfc_wire_236 (sink__dfc_wire_4821__dfc_wire_4799)
  );
  const_0x1_0000000000002000 const2045 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2153:90
    .clock                              (clock),
    .reset                              (reset),
    .const_fix_32_0_1__0000000000002000 (_const2045_const_fix_32_0_1__0000000000002000)
  );
  const_0x1_0000000000000620 const2060 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2154:90
    .clock                              (clock),
    .reset                              (reset),
    .const_fix_32_0_1__0000000000000620 (_const2060_const_fix_32_0_1__0000000000000620)
  );
  const_0x1_000000000000031f const2065 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2155:90
    .clock                              (clock),
    .reset                              (reset),
    .const_fix_32_0_1__000000000000031f (_const2065_const_fix_32_0_1__000000000000031f)
  );
  const_0x1_0000000000000fb1 const2068 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2156:90
    .clock                              (clock),
    .reset                              (reset),
    .const_fix_32_0_1__0000000000000fb1 (_const2068_const_fix_32_0_1__0000000000000fb1)
  );
  const_0x1_00000000000008e4 const2074 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2157:90
    .clock                              (clock),
    .reset                              (reset),
    .const_fix_32_0_1__00000000000008e4 (_const2074_const_fix_32_0_1__00000000000008e4)
  );
  const_0x1_0000000000000d4e const2081 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2158:90
    .clock                              (clock),
    .reset                              (reset),
    .const_fix_32_0_1__0000000000000d4e (_const2081_const_fix_32_0_1__0000000000000d4e)
  );
  const_0x1_ffffffffffffff00 const2086 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2159:90
    .clock                              (clock),
    .reset                              (reset),
    .const_fix_32_0_1__ffffffffffffff00 (_const2086_const_fix_32_0_1__ffffffffffffff00)
  );
  const_0x1_0000000000000968 const2097 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2160:90
    .clock                              (clock),
    .reset                              (reset),
    .const_fix_32_0_1__0000000000000968 (_const2097_const_fix_32_0_1__0000000000000968)
  );
  const_0x1_0000000000000ec8 const2098 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2161:90
    .clock                              (clock),
    .reset                              (reset),
    .const_fix_32_0_1__0000000000000ec8 (_const2098_const_fix_32_0_1__0000000000000ec8)
  );
  const_0x1_00000000000000b5 const2102 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2162:90
    .clock                              (clock),
    .reset                              (reset),
    .const_fix_32_0_1__00000000000000b5 (_const2102_const_fix_32_0_1__00000000000000b5)
  );
  const_0x1_0000000000000080 const2106 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2163:90
    .clock                              (clock),
    .reset                              (reset),
    .const_fix_32_0_1__0000000000000080 (_const2106_const_fix_32_0_1__0000000000000080)
  );
  const_0x1_0000000000000454 const2111 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2164:90
    .clock                              (clock),
    .reset                              (reset),
    .const_fix_32_0_1__0000000000000454 (_const2111_const_fix_32_0_1__0000000000000454)
  );
  const_0x1_0000000000000004 const2144 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2165:90
    .clock                              (clock),
    .reset                              (reset),
    .const_fix_32_0_1__0000000000000004 (_const2144_const_fix_32_0_1__0000000000000004)
  );
  const_0x1_00000000000000ff const2146 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2166:90
    .clock                              (clock),
    .reset                              (reset),
    .const_fix_32_0_1__00000000000000ff (_const2146_const_fix_32_0_1__00000000000000ff)
  );
  const_0x1_0000000000000235 const2149 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2167:90
    .clock                              (clock),
    .reset                              (reset),
    .const_fix_32_0_1__0000000000000235 (_const2149_const_fix_32_0_1__0000000000000235)
  );
  delay_fixed_32_0_1_996 delay_fixed_32_0_1_996_2150 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2168:146
    .clock (clock),
    .reset (reset),
    .in    (_dup49_const_fix_32_0_1__0000000000000235_4140),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
    .out   (_delay_fixed_32_0_1_996_2150_out)
  );
  delay_fixed_32_0_1_273 delay_fixed_32_0_1_273_2151 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2169:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1753__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1899:136
    .out   (_delay_fixed_32_0_1_273_2151_out)
  );
  delay_fixed_32_0_1_784 delay_fixed_32_0_1_784_2152 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2170:146
    .clock (clock),
    .reset (reset),
    .in    (_dup45_const_fix_32_0_1__0000000000000235_4140),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
    .out   (_delay_fixed_32_0_1_784_2152_out)
  );
  delay_fixed_32_0_1_917 delay_fixed_32_0_1_917_2153 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2171:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_4208),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_917_2153_out)
  );
  delay_fixed_32_0_1_962 delay_fixed_32_0_1_962_2154 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2172:146
    .clock (clock),
    .reset (reset),
    .in    (_dup43_const_fix_32_0_1__0000000000000235_4140),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
    .out   (_delay_fixed_32_0_1_962_2154_out)
  );
  delay_fixed_32_0_1_156 delay_fixed_32_0_1_156_2155 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2173:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1749__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1895:116
    .out   (_delay_fixed_32_0_1_156_2155_out)
  );
  delay_fixed_32_0_1_16 delay_fixed_32_0_1_16_2156 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2174:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1745__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1891:116
    .out   (_delay_fixed_32_0_1_16_2156_out)
  );
  delay_fixed_32_0_1_16 delay_fixed_32_0_1_16_2157 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2175:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1745__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1891:116
    .out   (_delay_fixed_32_0_1_16_2157_out)
  );
  delay_fixed_32_0_1_147 delay_fixed_32_0_1_147_2158 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2176:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1741__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1887:136
    .out   (_delay_fixed_32_0_1_147_2158_out)
  );
  delay_fixed_32_0_1_980 delay_fixed_32_0_1_980_2159 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2177:146
    .clock (clock),
    .reset (reset),
    .in    (_dup33_const_fix_32_0_1__0000000000000235_4140),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
    .out   (_delay_fixed_32_0_1_980_2159_out)
  );
  delay_fixed_32_0_1_240 delay_fixed_32_0_1_240_2160 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2178:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1737__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1883:136
    .out   (_delay_fixed_32_0_1_240_2160_out)
  );
  delay_fixed_32_0_1_876 delay_fixed_32_0_1_876_2161 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2179:146
    .clock (clock),
    .reset (reset),
    .in    (_dup29_const_fix_32_0_1__0000000000000235_4140),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
    .out   (_delay_fixed_32_0_1_876_2161_out)
  );
  delay_fixed_32_0_1_1007 delay_fixed_32_0_1_1007_2162 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2180:150
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_4172),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_1007_2162_out)
  );
  delay_fixed_32_0_1_1041 delay_fixed_32_0_1_1041_2163 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2181:150
    .clock (clock),
    .reset (reset),
    .in    (_dup27_const_fix_32_0_1__0000000000000235_4140),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
    .out   (_delay_fixed_32_0_1_1041_2163_out)
  );
  delay_fixed_32_0_1_46 delay_fixed_32_0_1_46_2164 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2182:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1732__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1878:116
    .out   (_delay_fixed_32_0_1_46_2164_out)
  );
  delay_fixed_32_0_1_436 delay_fixed_32_0_1_436_2165 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2183:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1729__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1875:136
    .out   (_delay_fixed_32_0_1_436_2165_out)
  );
  delay_fixed_32_0_1_825 delay_fixed_32_0_1_825_2166 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2184:146
    .clock (clock),
    .reset (reset),
    .in    (_dup21_const_fix_32_0_1__0000000000000235_4140),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
    .out   (_delay_fixed_32_0_1_825_2166_out)
  );
  delay_fixed_32_0_1_194 delay_fixed_32_0_1_194_2167 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2185:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1725__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1871:136
    .out   (_delay_fixed_32_0_1_194_2167_out)
  );
  delay_fixed_32_0_1_1055 delay_fixed_32_0_1_1055_2168 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2186:150
    .clock (clock),
    .reset (reset),
    .in    (_dup17_const_fix_32_0_1__0000000000000235_4140),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
    .out   (_delay_fixed_32_0_1_1055_2168_out)
  );
  delay_fixed_32_0_1_1099 delay_fixed_32_0_1_1099_2169 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2187:150
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_4144),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_1099_2169_out)
  );
  delay_fixed_32_0_1_1154 delay_fixed_32_0_1_1154_2170 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2188:150
    .clock (clock),
    .reset (reset),
    .in    (_dup15_const_fix_32_0_1__0000000000000235_4140),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
    .out   (_delay_fixed_32_0_1_1154_2170_out)
  );
  delay_fixed_32_0_1_274 delay_fixed_32_0_1_274_2171 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2189:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1721__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1867:116
    .out   (_delay_fixed_32_0_1_274_2171_out)
  );
  delay_fixed_32_0_1_990 delay_fixed_32_0_1_990_2172 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2190:146
    .clock (clock),
    .reset (reset),
    .in    (_dup821_const_fix_32_0_1__0000000000002000_4134),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:967:473
    .out   (_delay_fixed_32_0_1_990_2172_out)
  );
  delay_fixed_1_0_0_29 delay_fixed_1_0_0_29_2173 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2191:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1706__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1852:139
    .out   (_delay_fixed_1_0_0_29_2173_out)
  );
  delay_fixed_32_0_1_1596 delay_fixed_32_0_1_1596_2174 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2192:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4085),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1596_2174_out)
  );
  delay_fixed_32_0_1_1501 delay_fixed_32_0_1_1501_2175 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2193:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4081),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1501_2175_out)
  );
  delay_fixed_32_0_1_13 delay_fixed_32_0_1_13_2176 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2194:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1703__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1849:154
    .out   (_delay_fixed_32_0_1_13_2176_out)
  );
  delay_fixed_32_0_1_1548 delay_fixed_32_0_1_1548_2177 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2195:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4085),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1548_2177_out)
  );
  delay_fixed_32_0_1_1535 delay_fixed_32_0_1_1535_2178 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2196:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4081),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1535_2178_out)
  );
  delay_fixed_32_0_1_52 delay_fixed_32_0_1_52_2179 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2197:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1637__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1783:116
    .out   (_delay_fixed_32_0_1_52_2179_out)
  );
  delay_fixed_1_0_0_60 delay_fixed_1_0_0_60_2180 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2198:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1698__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1844:139
    .out   (_delay_fixed_1_0_0_60_2180_out)
  );
  delay_fixed_32_0_1_1812 delay_fixed_32_0_1_1812_2181 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2199:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4063),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1812_2181_out)
  );
  delay_fixed_32_0_1_1685 delay_fixed_32_0_1_1685_2182 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2200:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4059),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1685_2182_out)
  );
  delay_fixed_32_0_1_60 delay_fixed_32_0_1_60_2183 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2201:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1695__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1841:154
    .out   (_delay_fixed_32_0_1_60_2183_out)
  );
  delay_fixed_32_0_1_1779 delay_fixed_32_0_1_1779_2184 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2202:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4063),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1779_2184_out)
  );
  delay_fixed_32_0_1_1719 delay_fixed_32_0_1_1719_2185 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2203:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4059),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1719_2185_out)
  );
  delay_fixed_32_0_1_373 delay_fixed_32_0_1_373_2186 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2204:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1647__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1793:116
    .out   (_delay_fixed_32_0_1_373_2186_out)
  );
  delay_fixed_1_0_0_106 delay_fixed_1_0_0_106_2187 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2205:142
    .clock (clock),
    .reset (reset),
    .in    (_LT1690__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1836:139
    .out   (_delay_fixed_1_0_0_106_2187_out)
  );
  delay_fixed_32_0_1_1996 delay_fixed_32_0_1_1996_2188 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2206:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4041),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1996_2188_out)
  );
  delay_fixed_32_0_1_1831 delay_fixed_32_0_1_1831_2189 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2207:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4037),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1831_2189_out)
  );
  delay_fixed_32_0_1_75 delay_fixed_32_0_1_75_2190 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2208:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1687__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1833:154
    .out   (_delay_fixed_32_0_1_75_2190_out)
  );
  delay_fixed_32_0_1_1940 delay_fixed_32_0_1_1940_2191 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2209:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4041),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1940_2191_out)
  );
  delay_fixed_32_0_1_1865 delay_fixed_32_0_1_1865_2192 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2210:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4037),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1865_2192_out)
  );
  delay_fixed_32_0_1_388 delay_fixed_32_0_1_388_2193 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2211:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1657__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1803:116
    .out   (_delay_fixed_32_0_1_388_2193_out)
  );
  delay_fixed_32_0_1_29 delay_fixed_32_0_1_29_2194 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2212:142
    .clock (clock),
    .reset (reset),
    .in    (_MUX1681__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1827:169
    .out   (_delay_fixed_32_0_1_29_2194_out)
  );
  delay_fixed_32_0_1_1391 delay_fixed_32_0_1_1391_2195 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2213:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4019),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1391_2195_out)
  );
  delay_fixed_32_0_1_1337 delay_fixed_32_0_1_1337_2196 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2214:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4015),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1337_2196_out)
  );
  delay_fixed_32_0_1_20 delay_fixed_32_0_1_20_2197 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2215:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1679__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1825:154
    .out   (_delay_fixed_32_0_1_20_2197_out)
  );
  delay_fixed_32_0_1_1391 delay_fixed_32_0_1_1391_2198 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2216:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4019),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1391_2198_out)
  );
  delay_fixed_32_0_1_1371 delay_fixed_32_0_1_1371_2199 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2217:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4015),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1371_2199_out)
  );
  delay_fixed_32_0_1_84 delay_fixed_32_0_1_84_2200 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2218:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1667__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1813:116
    .out   (_delay_fixed_32_0_1_84_2200_out)
  );
  delay_fixed_32_0_1_26 delay_fixed_32_0_1_26_2201 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2219:142
    .clock (clock),
    .reset (reset),
    .in    (_MUX1673__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1819:169
    .out   (_delay_fixed_32_0_1_26_2201_out)
  );
  delay_fixed_32_0_1_1446 delay_fixed_32_0_1_1446_2202 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2220:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3997),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1446_2202_out)
  );
  delay_fixed_32_0_1_1407 delay_fixed_32_0_1_1407_2203 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2221:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3993),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1407_2203_out)
  );
  delay_fixed_32_0_1_11 delay_fixed_32_0_1_11_2204 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2222:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1671__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1817:154
    .out   (_delay_fixed_32_0_1_11_2204_out)
  );
  delay_fixed_32_0_1_1452 delay_fixed_32_0_1_1452_2205 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2223:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3997),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1452_2205_out)
  );
  delay_fixed_32_0_1_1441 delay_fixed_32_0_1_1441_2206 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2224:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3993),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1441_2206_out)
  );
  delay_fixed_32_0_1_84 delay_fixed_32_0_1_84_2207 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2225:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1667__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1813:116
    .out   (_delay_fixed_32_0_1_84_2207_out)
  );
  delay_fixed_1_0_0_86 delay_fixed_1_0_0_86_2208 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2226:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1664__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1810:139
    .out   (_delay_fixed_1_0_0_86_2208_out)
  );
  delay_fixed_32_0_1_1848 delay_fixed_32_0_1_1848_2209 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2227:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3975),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1848_2209_out)
  );
  delay_fixed_32_0_1_1729 delay_fixed_32_0_1_1729_2210 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2228:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3971),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1729_2210_out)
  );
  delay_fixed_32_0_1_41 delay_fixed_32_0_1_41_2211 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2229:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1661__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1807:154
    .out   (_delay_fixed_32_0_1_41_2211_out)
  );
  delay_fixed_32_0_1_1804 delay_fixed_32_0_1_1804_2212 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2230:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3975),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1804_2212_out)
  );
  delay_fixed_32_0_1_1763 delay_fixed_32_0_1_1763_2213 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2231:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3971),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1763_2213_out)
  );
  delay_fixed_32_0_1_388 delay_fixed_32_0_1_388_2214 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2232:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1657__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1803:116
    .out   (_delay_fixed_32_0_1_388_2214_out)
  );
  delay_fixed_1_0_0_5 delay_fixed_1_0_0_5_2215 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2233:134
    .clock (clock),
    .reset (reset),
    .in    (_LT1654__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1800:139
    .out   (_delay_fixed_1_0_0_5_2215_out)
  );
  delay_fixed_32_0_1_1790 delay_fixed_32_0_1_1790_2216 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2234:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3953),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1790_2216_out)
  );
  delay_fixed_32_0_1_1722 delay_fixed_32_0_1_1722_2217 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2235:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3949),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1722_2217_out)
  );
  delay_fixed_32_0_1_19 delay_fixed_32_0_1_19_2218 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2236:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1651__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1797:154
    .out   (_delay_fixed_32_0_1_19_2218_out)
  );
  delay_fixed_32_0_1_1775 delay_fixed_32_0_1_1775_2219 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2237:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3953),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1775_2219_out)
  );
  delay_fixed_32_0_1_1756 delay_fixed_32_0_1_1756_2220 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2238:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3949),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1756_2220_out)
  );
  delay_fixed_32_0_1_373 delay_fixed_32_0_1_373_2221 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2239:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1647__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1793:116
    .out   (_delay_fixed_32_0_1_373_2221_out)
  );
  delay_fixed_1_0_0_92 delay_fixed_1_0_0_92_2222 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2240:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1644__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1790:139
    .out   (_delay_fixed_1_0_0_92_2222_out)
  );
  delay_fixed_32_0_1_1612 delay_fixed_32_0_1_1612_2223 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2241:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3931),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1612_2223_out)
  );
  delay_fixed_32_0_1_1483 delay_fixed_32_0_1_1483_2224 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2242:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3927),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1483_2224_out)
  );
  delay_fixed_32_0_1_62 delay_fixed_32_0_1_62_2225 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2243:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1641__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1787:154
    .out   (_delay_fixed_32_0_1_62_2225_out)
  );
  delay_fixed_32_0_1_1579 delay_fixed_32_0_1_1579_2226 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2244:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3931),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1579_2226_out)
  );
  delay_fixed_32_0_1_1517 delay_fixed_32_0_1_1517_2227 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2245:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3927),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1517_2227_out)
  );
  delay_fixed_32_0_1_52 delay_fixed_32_0_1_52_2228 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2246:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1637__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1783:116
    .out   (_delay_fixed_32_0_1_52_2228_out)
  );
  delay_fixed_32_0_1_1561 delay_fixed_32_0_1_1561_2229 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2247:150
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_3916),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_1561_2229_out)
  );
  delay_fixed_32_0_1_1421 delay_fixed_32_0_1_1421_2230 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2248:150
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_3912),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_1421_2230_out)
  );
  delay_fixed_32_0_1_21 delay_fixed_32_0_1_21_2231 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2249:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1627__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1773:116
    .out   (_delay_fixed_32_0_1_21_2231_out)
  );
  delay_fixed_32_0_1_1478 delay_fixed_32_0_1_1478_2232 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2250:150
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_3904),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_1478_2232_out)
  );
  delay_fixed_32_0_1_1365 delay_fixed_32_0_1_1365_2233 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2251:150
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_3900),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_1365_2233_out)
  );
  delay_fixed_32_0_1_21 delay_fixed_32_0_1_21_2234 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2252:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1627__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1773:116
    .out   (_delay_fixed_32_0_1_21_2234_out)
  );
  delay_fixed_32_0_1_102 delay_fixed_32_0_1_102_2235 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2253:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1623__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1769:116
    .out   (_delay_fixed_32_0_1_102_2235_out)
  );
  delay_fixed_32_0_1_102 delay_fixed_32_0_1_102_2236 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2254:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1623__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1769:116
    .out   (_delay_fixed_32_0_1_102_2236_out)
  );
  delay_fixed_32_0_1_65 delay_fixed_32_0_1_65_2237 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2255:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1619__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1765:116
    .out   (_delay_fixed_32_0_1_65_2237_out)
  );
  delay_fixed_32_0_1_65 delay_fixed_32_0_1_65_2238 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2256:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1619__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1765:116
    .out   (_delay_fixed_32_0_1_65_2238_out)
  );
  delay_fixed_32_0_1_71 delay_fixed_32_0_1_71_2239 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2257:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1616__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1762:116
    .out   (_delay_fixed_32_0_1_71_2239_out)
  );
  delay_fixed_32_0_1_71 delay_fixed_32_0_1_71_2240 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2258:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1616__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1762:116
    .out   (_delay_fixed_32_0_1_71_2240_out)
  );
  delay_fixed_32_0_1_145 delay_fixed_32_0_1_145_2241 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2259:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1612__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1758:116
    .out   (_delay_fixed_32_0_1_145_2241_out)
  );
  delay_fixed_32_0_1_145 delay_fixed_32_0_1_145_2242 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2260:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1612__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1758:116
    .out   (_delay_fixed_32_0_1_145_2242_out)
  );
  delay_fixed_32_0_1_17 delay_fixed_32_0_1_17_2243 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2261:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL1608__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1754:136
    .out   (_delay_fixed_32_0_1_17_2243_out)
  );
  delay_fixed_32_0_1_1013 delay_fixed_32_0_1_1013_2244 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2262:150
    .clock (clock),
    .reset (reset),
    .in    (_dup49_const_fix_32_0_1__0000000000000235_3776),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
    .out   (_delay_fixed_32_0_1_1013_2244_out)
  );
  delay_fixed_32_0_1_114 delay_fixed_32_0_1_114_2245 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2263:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1604__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1750:136
    .out   (_delay_fixed_32_0_1_114_2245_out)
  );
  delay_fixed_32_0_1_871 delay_fixed_32_0_1_871_2246 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2264:146
    .clock (clock),
    .reset (reset),
    .in    (_dup45_const_fix_32_0_1__0000000000000235_3776),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
    .out   (_delay_fixed_32_0_1_871_2246_out)
  );
  delay_fixed_32_0_1_898 delay_fixed_32_0_1_898_2247 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2265:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_3844),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_898_2247_out)
  );
  delay_fixed_32_0_1_986 delay_fixed_32_0_1_986_2248 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2266:146
    .clock (clock),
    .reset (reset),
    .in    (_dup43_const_fix_32_0_1__0000000000000235_3776),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
    .out   (_delay_fixed_32_0_1_986_2248_out)
  );
  delay_fixed_32_0_1_86 delay_fixed_32_0_1_86_2249 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2267:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1600__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1746:116
    .out   (_delay_fixed_32_0_1_86_2249_out)
  );
  delay_fixed_32_0_1_7 delay_fixed_32_0_1_7_2250 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2268:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1596__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1742:116
    .out   (_delay_fixed_32_0_1_7_2250_out)
  );
  delay_fixed_32_0_1_7 delay_fixed_32_0_1_7_2251 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2269:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1596__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1742:116
    .out   (_delay_fixed_32_0_1_7_2251_out)
  );
  delay_fixed_32_0_1_71 delay_fixed_32_0_1_71_2252 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2270:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL1592__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1738:136
    .out   (_delay_fixed_32_0_1_71_2252_out)
  );
  delay_fixed_32_0_1_906 delay_fixed_32_0_1_906_2253 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2271:146
    .clock (clock),
    .reset (reset),
    .in    (_dup33_const_fix_32_0_1__0000000000000235_3776),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
    .out   (_delay_fixed_32_0_1_906_2253_out)
  );
  delay_fixed_32_0_1_67 delay_fixed_32_0_1_67_2254 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2272:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL1588__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1734:136
    .out   (_delay_fixed_32_0_1_67_2254_out)
  );
  delay_fixed_32_0_1_819 delay_fixed_32_0_1_819_2255 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2273:146
    .clock (clock),
    .reset (reset),
    .in    (_dup29_const_fix_32_0_1__0000000000000235_3776),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
    .out   (_delay_fixed_32_0_1_819_2255_out)
  );
  delay_fixed_32_0_1_908 delay_fixed_32_0_1_908_2256 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2274:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_3808),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_908_2256_out)
  );
  delay_fixed_32_0_1_965 delay_fixed_32_0_1_965_2257 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2275:146
    .clock (clock),
    .reset (reset),
    .in    (_dup27_const_fix_32_0_1__0000000000000235_3776),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
    .out   (_delay_fixed_32_0_1_965_2257_out)
  );
  delay_fixed_32_0_1_29 delay_fixed_32_0_1_29_2258 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2276:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1583__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1729:116
    .out   (_delay_fixed_32_0_1_29_2258_out)
  );
  delay_fixed_32_0_1_130 delay_fixed_32_0_1_130_2259 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2277:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1580__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1726:136
    .out   (_delay_fixed_32_0_1_130_2259_out)
  );
  delay_fixed_32_0_1_913 delay_fixed_32_0_1_913_2260 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2278:146
    .clock (clock),
    .reset (reset),
    .in    (_dup21_const_fix_32_0_1__0000000000000235_3776),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
    .out   (_delay_fixed_32_0_1_913_2260_out)
  );
  delay_fixed_32_0_1_155 delay_fixed_32_0_1_155_2261 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2279:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1576__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1722:136
    .out   (_delay_fixed_32_0_1_155_2261_out)
  );
  delay_fixed_32_0_1_837 delay_fixed_32_0_1_837_2262 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2280:146
    .clock (clock),
    .reset (reset),
    .in    (_dup17_const_fix_32_0_1__0000000000000235_3776),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
    .out   (_delay_fixed_32_0_1_837_2262_out)
  );
  delay_fixed_32_0_1_838 delay_fixed_32_0_1_838_2263 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2281:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_3780),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_838_2263_out)
  );
  delay_fixed_32_0_1_886 delay_fixed_32_0_1_886_2264 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2282:146
    .clock (clock),
    .reset (reset),
    .in    (_dup15_const_fix_32_0_1__0000000000000235_3776),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
    .out   (_delay_fixed_32_0_1_886_2264_out)
  );
  delay_fixed_32_0_1_32 delay_fixed_32_0_1_32_2265 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2283:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1571__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1717:116
    .out   (_delay_fixed_32_0_1_32_2265_out)
  );
  delay_fixed_32_0_1_923 delay_fixed_32_0_1_923_2266 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2284:146
    .clock (clock),
    .reset (reset),
    .in    (_dup821_const_fix_32_0_1__0000000000002000_3770),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:967:473
    .out   (_delay_fixed_32_0_1_923_2266_out)
  );
  delay_fixed_1_0_0_42 delay_fixed_1_0_0_42_2267 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2285:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1557__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1703:139
    .out   (_delay_fixed_1_0_0_42_2267_out)
  );
  delay_fixed_32_0_1_1392 delay_fixed_32_0_1_1392_2268 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2286:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3721),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1392_2268_out)
  );
  delay_fixed_32_0_1_1304 delay_fixed_32_0_1_1304_2269 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2287:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3717),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1304_2269_out)
  );
  delay_fixed_32_0_1_31 delay_fixed_32_0_1_31_2270 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2288:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1554__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1700:154
    .out   (_delay_fixed_32_0_1_31_2270_out)
  );
  delay_fixed_32_0_1_1369 delay_fixed_32_0_1_1369_2271 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2289:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3721),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1369_2271_out)
  );
  delay_fixed_32_0_1_1338 delay_fixed_32_0_1_1338_2272 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2290:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3717),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1338_2272_out)
  );
  delay_fixed_32_0_1_6 delay_fixed_32_0_1_6_2273 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2291:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1488__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1634:116
    .out   (_delay_fixed_32_0_1_6_2273_out)
  );
  delay_fixed_1_0_0_114 delay_fixed_1_0_0_114_2274 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2292:142
    .clock (clock),
    .reset (reset),
    .in    (_LT1549__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1695:139
    .out   (_delay_fixed_1_0_0_114_2274_out)
  );
  delay_fixed_32_0_1_1771 delay_fixed_32_0_1_1771_2275 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2293:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3699),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1771_2275_out)
  );
  delay_fixed_32_0_1_1632 delay_fixed_32_0_1_1632_2276 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2294:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3695),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1632_2276_out)
  );
  delay_fixed_32_0_1_75 delay_fixed_32_0_1_75_2277 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2295:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1546__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1692:154
    .out   (_delay_fixed_32_0_1_75_2277_out)
  );
  delay_fixed_32_0_1_1741 delay_fixed_32_0_1_1741_2278 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2296:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3699),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1741_2278_out)
  );
  delay_fixed_32_0_1_1666 delay_fixed_32_0_1_1666_2279 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2297:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3695),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1666_2279_out)
  );
  delay_fixed_32_0_1_248 delay_fixed_32_0_1_248_2280 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2298:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1498__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1644:116
    .out   (_delay_fixed_32_0_1_248_2280_out)
  );
  delay_fixed_1_0_0_25 delay_fixed_1_0_0_25_2281 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2299:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1541__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1687:139
    .out   (_delay_fixed_1_0_0_25_2281_out)
  );
  delay_fixed_32_0_1_1691 delay_fixed_32_0_1_1691_2282 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2300:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3677),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1691_2282_out)
  );
  delay_fixed_32_0_1_1628 delay_fixed_32_0_1_1628_2283 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2301:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3673),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1628_2283_out)
  );
  delay_fixed_32_0_1_13 delay_fixed_32_0_1_13_2284 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2302:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1538__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1684:154
    .out   (_delay_fixed_32_0_1_13_2284_out)
  );
  delay_fixed_32_0_1_1675 delay_fixed_32_0_1_1675_2285 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2303:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3677),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1675_2285_out)
  );
  delay_fixed_32_0_1_1662 delay_fixed_32_0_1_1662_2286 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2304:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3673),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1662_2286_out)
  );
  delay_fixed_32_0_1_26 delay_fixed_32_0_1_26_2287 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2305:142
    .clock (clock),
    .reset (reset),
    .in    (_MUX1524__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1670:169
    .out   (_delay_fixed_32_0_1_26_2287_out)
  );
  delay_fixed_32_0_1_1449 delay_fixed_32_0_1_1449_2288 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2306:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3633),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1449_2288_out)
  );
  delay_fixed_32_0_1_1368 delay_fixed_32_0_1_1368_2289 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2307:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3629),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1368_2289_out)
  );
  delay_fixed_32_0_1_6 delay_fixed_32_0_1_6_2290 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2308:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1522__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1668:154
    .out   (_delay_fixed_32_0_1_6_2290_out)
  );
  delay_fixed_32_0_1_1408 delay_fixed_32_0_1_1408_2291 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2309:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3633),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1408_2291_out)
  );
  delay_fixed_32_0_1_1402 delay_fixed_32_0_1_1402_2292 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2310:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3629),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1402_2292_out)
  );
  delay_fixed_32_0_1_23 delay_fixed_32_0_1_23_2293 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2311:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1518__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1664:116
    .out   (_delay_fixed_32_0_1_23_2293_out)
  );
  delay_fixed_32_0_1_1643 delay_fixed_32_0_1_1643_2294 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2312:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3585),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1643_2294_out)
  );
  delay_fixed_32_0_1_248 delay_fixed_32_0_1_248_2295 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2313:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1498__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1644:116
    .out   (_delay_fixed_32_0_1_248_2295_out)
  );
  delay_fixed_1_0_0_63 delay_fixed_1_0_0_63_2296 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2314:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1495__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1641:139
    .out   (_delay_fixed_1_0_0_63_2296_out)
  );
  delay_fixed_32_0_1_1341 delay_fixed_32_0_1_1341_2297 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2315:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3567),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1341_2297_out)
  );
  delay_fixed_32_0_1_1267 delay_fixed_32_0_1_1267_2298 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2316:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3563),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1267_2298_out)
  );
  delay_fixed_32_0_1_53 delay_fixed_32_0_1_53_2299 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2317:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1492__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1638:154
    .out   (_delay_fixed_32_0_1_53_2299_out)
  );
  delay_fixed_32_0_1_1354 delay_fixed_32_0_1_1354_2300 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2318:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3567),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1354_2300_out)
  );
  delay_fixed_32_0_1_1301 delay_fixed_32_0_1_1301_2301 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2319:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3563),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1301_2301_out)
  );
  delay_fixed_32_0_1_6 delay_fixed_32_0_1_6_2302 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2320:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1488__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1634:116
    .out   (_delay_fixed_32_0_1_6_2302_out)
  );
  delay_fixed_32_0_1_1488 delay_fixed_32_0_1_1488_2303 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2321:150
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_3552),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_1488_2303_out)
  );
  delay_fixed_32_0_1_1323 delay_fixed_32_0_1_1323_2304 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2322:150
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_3548),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_1323_2304_out)
  );
  delay_fixed_32_0_1_172 delay_fixed_32_0_1_172_2305 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2323:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1478__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1624:116
    .out   (_delay_fixed_32_0_1_172_2305_out)
  );
  delay_fixed_32_0_1_1391 delay_fixed_32_0_1_1391_2306 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2324:150
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_3540),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_1391_2306_out)
  );
  delay_fixed_32_0_1_1316 delay_fixed_32_0_1_1316_2307 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2325:150
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_3536),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_1316_2307_out)
  );
  delay_fixed_32_0_1_172 delay_fixed_32_0_1_172_2308 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2326:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1478__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1624:116
    .out   (_delay_fixed_32_0_1_172_2308_out)
  );
  delay_fixed_32_0_1_49 delay_fixed_32_0_1_49_2309 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2327:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1474__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1620:116
    .out   (_delay_fixed_32_0_1_49_2309_out)
  );
  delay_fixed_32_0_1_49 delay_fixed_32_0_1_49_2310 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2328:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1474__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1620:116
    .out   (_delay_fixed_32_0_1_49_2310_out)
  );
  delay_fixed_32_0_1_119 delay_fixed_32_0_1_119_2311 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2329:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1470__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1616:116
    .out   (_delay_fixed_32_0_1_119_2311_out)
  );
  delay_fixed_32_0_1_119 delay_fixed_32_0_1_119_2312 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2330:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1470__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1616:116
    .out   (_delay_fixed_32_0_1_119_2312_out)
  );
  delay_fixed_32_0_1_27 delay_fixed_32_0_1_27_2313 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2331:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1466__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1612:116
    .out   (_delay_fixed_32_0_1_27_2313_out)
  );
  delay_fixed_32_0_1_27 delay_fixed_32_0_1_27_2314 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2332:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1466__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1612:116
    .out   (_delay_fixed_32_0_1_27_2314_out)
  );
  delay_fixed_32_0_1_11 delay_fixed_32_0_1_11_2315 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2333:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1463__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1609:116
    .out   (_delay_fixed_32_0_1_11_2315_out)
  );
  delay_fixed_32_0_1_11 delay_fixed_32_0_1_11_2316 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2334:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1463__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1609:116
    .out   (_delay_fixed_32_0_1_11_2316_out)
  );
  delay_fixed_32_0_1_109 delay_fixed_32_0_1_109_2317 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2335:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1459__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1605:136
    .out   (_delay_fixed_32_0_1_109_2317_out)
  );
  delay_fixed_32_0_1_853 delay_fixed_32_0_1_853_2318 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2336:146
    .clock (clock),
    .reset (reset),
    .in    (_dup49_const_fix_32_0_1__0000000000000235_3412),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
    .out   (_delay_fixed_32_0_1_853_2318_out)
  );
  delay_fixed_32_0_1_274 delay_fixed_32_0_1_274_2319 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2337:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1455__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1601:136
    .out   (_delay_fixed_32_0_1_274_2319_out)
  );
  delay_fixed_32_0_1_644 delay_fixed_32_0_1_644_2320 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2338:146
    .clock (clock),
    .reset (reset),
    .in    (_dup45_const_fix_32_0_1__0000000000000235_3412),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
    .out   (_delay_fixed_32_0_1_644_2320_out)
  );
  delay_fixed_32_0_1_732 delay_fixed_32_0_1_732_2321 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2339:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_3480),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_732_2321_out)
  );
  delay_fixed_32_0_1_825 delay_fixed_32_0_1_825_2322 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2340:146
    .clock (clock),
    .reset (reset),
    .in    (_dup43_const_fix_32_0_1__0000000000000235_3412),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
    .out   (_delay_fixed_32_0_1_825_2322_out)
  );
  delay_fixed_32_0_1_153 delay_fixed_32_0_1_153_2323 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2341:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1451__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1597:116
    .out   (_delay_fixed_32_0_1_153_2323_out)
  );
  delay_fixed_32_0_1_160 delay_fixed_32_0_1_160_2324 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2342:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1447__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1593:116
    .out   (_delay_fixed_32_0_1_160_2324_out)
  );
  delay_fixed_32_0_1_160 delay_fixed_32_0_1_160_2325 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2343:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1447__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1593:116
    .out   (_delay_fixed_32_0_1_160_2325_out)
  );
  delay_fixed_32_0_1_171 delay_fixed_32_0_1_171_2326 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2344:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1443__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1589:136
    .out   (_delay_fixed_32_0_1_171_2326_out)
  );
  delay_fixed_32_0_1_681 delay_fixed_32_0_1_681_2327 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2345:146
    .clock (clock),
    .reset (reset),
    .in    (_dup33_const_fix_32_0_1__0000000000000235_3412),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
    .out   (_delay_fixed_32_0_1_681_2327_out)
  );
  delay_fixed_32_0_1_92 delay_fixed_32_0_1_92_2328 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2346:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL1439__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1585:136
    .out   (_delay_fixed_32_0_1_92_2328_out)
  );
  delay_fixed_32_0_1_668 delay_fixed_32_0_1_668_2329 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2347:146
    .clock (clock),
    .reset (reset),
    .in    (_dup29_const_fix_32_0_1__0000000000000235_3412),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
    .out   (_delay_fixed_32_0_1_668_2329_out)
  );
  delay_fixed_32_0_1_666 delay_fixed_32_0_1_666_2330 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2348:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_3444),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_666_2330_out)
  );
  delay_fixed_32_0_1_779 delay_fixed_32_0_1_779_2331 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2349:146
    .clock (clock),
    .reset (reset),
    .in    (_dup27_const_fix_32_0_1__0000000000000235_3412),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
    .out   (_delay_fixed_32_0_1_779_2331_out)
  );
  delay_fixed_32_0_1_45 delay_fixed_32_0_1_45_2332 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2350:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1435__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1581:116
    .out   (_delay_fixed_32_0_1_45_2332_out)
  );
  delay_fixed_32_0_1_163 delay_fixed_32_0_1_163_2333 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2351:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1431__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1577:136
    .out   (_delay_fixed_32_0_1_163_2333_out)
  );
  delay_fixed_32_0_1_765 delay_fixed_32_0_1_765_2334 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2352:146
    .clock (clock),
    .reset (reset),
    .in    (_dup21_const_fix_32_0_1__0000000000000235_3412),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
    .out   (_delay_fixed_32_0_1_765_2334_out)
  );
  delay_fixed_32_0_1_152 delay_fixed_32_0_1_152_2335 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2353:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1427__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1573:136
    .out   (_delay_fixed_32_0_1_152_2335_out)
  );
  delay_fixed_32_0_1_708 delay_fixed_32_0_1_708_2336 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2354:146
    .clock (clock),
    .reset (reset),
    .in    (_dup17_const_fix_32_0_1__0000000000000235_3412),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
    .out   (_delay_fixed_32_0_1_708_2336_out)
  );
  delay_fixed_32_0_1_778 delay_fixed_32_0_1_778_2337 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2355:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_3416),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_778_2337_out)
  );
  delay_fixed_32_0_1_772 delay_fixed_32_0_1_772_2338 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2356:146
    .clock (clock),
    .reset (reset),
    .in    (_dup15_const_fix_32_0_1__0000000000000235_3412),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
    .out   (_delay_fixed_32_0_1_772_2338_out)
  );
  delay_fixed_32_0_1_13 delay_fixed_32_0_1_13_2339 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2357:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1422__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1568:116
    .out   (_delay_fixed_32_0_1_13_2339_out)
  );
  delay_fixed_32_0_1_902 delay_fixed_32_0_1_902_2340 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2358:146
    .clock (clock),
    .reset (reset),
    .in    (_dup821_const_fix_32_0_1__0000000000002000_3406),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:967:473
    .out   (_delay_fixed_32_0_1_902_2340_out)
  );
  delay_fixed_1_0_0_55 delay_fixed_1_0_0_55_2341 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2359:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1408__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1554:139
    .out   (_delay_fixed_1_0_0_55_2341_out)
  );
  delay_fixed_32_0_1_1306 delay_fixed_32_0_1_1306_2342 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2360:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3357),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1306_2342_out)
  );
  delay_fixed_32_0_1_1234 delay_fixed_32_0_1_1234_2343 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2361:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3353),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1234_2343_out)
  );
  delay_fixed_32_0_1_52 delay_fixed_32_0_1_52_2344 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2362:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1405__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1551:154
    .out   (_delay_fixed_32_0_1_52_2344_out)
  );
  delay_fixed_32_0_1_1320 delay_fixed_32_0_1_1320_2345 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2363:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3357),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1320_2345_out)
  );
  delay_fixed_32_0_1_1268 delay_fixed_32_0_1_1268_2346 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2364:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3353),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1268_2346_out)
  );
  delay_fixed_32_0_1_48 delay_fixed_32_0_1_48_2347 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2365:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1340__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1486:116
    .out   (_delay_fixed_32_0_1_48_2347_out)
  );
  delay_fixed_1_0_0_43 delay_fixed_1_0_0_43_2348 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2366:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1400__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1546:139
    .out   (_delay_fixed_1_0_0_43_2348_out)
  );
  delay_fixed_32_0_1_1626 delay_fixed_32_0_1_1626_2349 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2367:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3335),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1626_2349_out)
  );
  delay_fixed_32_0_1_1523 delay_fixed_32_0_1_1523_2350 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2368:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3331),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1523_2350_out)
  );
  delay_fixed_32_0_1_45 delay_fixed_32_0_1_45_2351 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2369:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1397__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1543:154
    .out   (_delay_fixed_32_0_1_45_2351_out)
  );
  delay_fixed_32_0_1_1602 delay_fixed_32_0_1_1602_2352 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2370:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3335),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1602_2352_out)
  );
  delay_fixed_32_0_1_1557 delay_fixed_32_0_1_1557_2353 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2371:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3331),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1557_2353_out)
  );
  delay_fixed_32_0_1_59 delay_fixed_32_0_1_59_2354 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2372:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1349__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1495:116
    .out   (_delay_fixed_32_0_1_59_2354_out)
  );
  delay_fixed_1_0_0_48 delay_fixed_1_0_0_48_2355 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2373:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1392__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1538:139
    .out   (_delay_fixed_1_0_0_48_2355_out)
  );
  delay_fixed_32_0_1_1604 delay_fixed_32_0_1_1604_2356 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2374:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3313),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1604_2356_out)
  );
  delay_fixed_32_0_1_1486 delay_fixed_32_0_1_1486_2357 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2375:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3309),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1486_2357_out)
  );
  delay_fixed_32_0_1_35 delay_fixed_32_0_1_35_2358 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2376:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1389__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1535:154
    .out   (_delay_fixed_32_0_1_35_2358_out)
  );
  delay_fixed_32_0_1_1555 delay_fixed_32_0_1_1555_2359 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2377:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3313),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1555_2359_out)
  );
  delay_fixed_32_0_1_1520 delay_fixed_32_0_1_1520_2360 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2378:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3309),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1520_2360_out)
  );
  delay_fixed_32_0_1_18 delay_fixed_32_0_1_18_2361 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2379:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1359__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1505:116
    .out   (_delay_fixed_32_0_1_18_2361_out)
  );
  delay_fixed_1_0_0_71 delay_fixed_1_0_0_71_2362 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2380:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1384__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1530:139
    .out   (_delay_fixed_1_0_0_71_2362_out)
  );
  delay_fixed_32_0_1_1487 delay_fixed_32_0_1_1487_2363 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2381:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3291),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1487_2363_out)
  );
  delay_fixed_32_0_1_1360 delay_fixed_32_0_1_1360_2364 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2382:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3287),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1360_2364_out)
  );
  delay_fixed_32_0_1_55 delay_fixed_32_0_1_55_2365 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2383:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1381__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1527:154
    .out   (_delay_fixed_32_0_1_55_2365_out)
  );
  delay_fixed_32_0_1_1449 delay_fixed_32_0_1_1449_2366 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2384:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3291),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1449_2366_out)
  );
  delay_fixed_32_0_1_1394 delay_fixed_32_0_1_1394_2367 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2385:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3287),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1394_2367_out)
  );
  delay_fixed_32_0_1_159 delay_fixed_32_0_1_159_2368 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2386:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1370__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1516:116
    .out   (_delay_fixed_32_0_1_159_2368_out)
  );
  delay_fixed_1_0_0_114 delay_fixed_1_0_0_114_2369 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2387:142
    .clock (clock),
    .reset (reset),
    .in    (_LT1376__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1522:139
    .out   (_delay_fixed_1_0_0_114_2369_out)
  );
  delay_fixed_32_0_1_1450 delay_fixed_32_0_1_1450_2370 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2388:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3269),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1450_2370_out)
  );
  delay_fixed_32_0_1_1326 delay_fixed_32_0_1_1326_2371 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2389:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3265),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1326_2371_out)
  );
  delay_fixed_32_0_1_31 delay_fixed_32_0_1_31_2372 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2390:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1373__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1519:154
    .out   (_delay_fixed_32_0_1_31_2372_out)
  );
  delay_fixed_32_0_1_1391 delay_fixed_32_0_1_1391_2373 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2391:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3269),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1391_2373_out)
  );
  delay_fixed_32_0_1_1360 delay_fixed_32_0_1_1360_2374 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2392:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3265),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1360_2374_out)
  );
  delay_fixed_32_0_1_159 delay_fixed_32_0_1_159_2375 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2393:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1370__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1516:116
    .out   (_delay_fixed_32_0_1_159_2375_out)
  );
  delay_fixed_1_0_0_64 delay_fixed_1_0_0_64_2376 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2394:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1366__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1512:139
    .out   (_delay_fixed_1_0_0_64_2376_out)
  );
  delay_fixed_32_0_1_1540 delay_fixed_32_0_1_1540_2377 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2395:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3247),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1540_2377_out)
  );
  delay_fixed_32_0_1_1429 delay_fixed_32_0_1_1429_2378 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2396:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3243),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1429_2378_out)
  );
  delay_fixed_32_0_1_56 delay_fixed_32_0_1_56_2379 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2397:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1363__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1509:154
    .out   (_delay_fixed_32_0_1_56_2379_out)
  );
  delay_fixed_32_0_1_1519 delay_fixed_32_0_1_1519_2380 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2398:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3247),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1519_2380_out)
  );
  delay_fixed_32_0_1_1463 delay_fixed_32_0_1_1463_2381 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2399:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3243),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1463_2381_out)
  );
  delay_fixed_32_0_1_18 delay_fixed_32_0_1_18_2382 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2400:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1359__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1505:116
    .out   (_delay_fixed_32_0_1_18_2382_out)
  );
  delay_fixed_1_0_0_101 delay_fixed_1_0_0_101_2383 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2401:142
    .clock (clock),
    .reset (reset),
    .in    (_LT1356__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1502:139
    .out   (_delay_fixed_1_0_0_101_2383_out)
  );
  delay_fixed_32_0_1_1602 delay_fixed_32_0_1_1602_2384 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2402:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3225),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1602_2384_out)
  );
  delay_fixed_32_0_1_1462 delay_fixed_32_0_1_1462_2385 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2403:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3221),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1462_2385_out)
  );
  delay_fixed_32_0_1_55 delay_fixed_32_0_1_55_2386 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2404:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1353__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1499:154
    .out   (_delay_fixed_32_0_1_55_2386_out)
  );
  delay_fixed_32_0_1_1551 delay_fixed_32_0_1_1551_2387 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2405:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3225),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1551_2387_out)
  );
  delay_fixed_32_0_1_1496 delay_fixed_32_0_1_1496_2388 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2406:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3221),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1496_2388_out)
  );
  delay_fixed_32_0_1_59 delay_fixed_32_0_1_59_2389 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2407:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1349__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1495:116
    .out   (_delay_fixed_32_0_1_59_2389_out)
  );
  delay_fixed_1_0_0_101 delay_fixed_1_0_0_101_2390 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2408:142
    .clock (clock),
    .reset (reset),
    .in    (_LT1346__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1492:139
    .out   (_delay_fixed_1_0_0_101_2390_out)
  );
  delay_fixed_32_0_1_1410 delay_fixed_32_0_1_1410_2391 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2409:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3203),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1410_2391_out)
  );
  delay_fixed_32_0_1_1227 delay_fixed_32_0_1_1227_2392 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2410:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3199),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1227_2392_out)
  );
  delay_fixed_32_0_1_96 delay_fixed_32_0_1_96_2393 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2411:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1343__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1489:154
    .out   (_delay_fixed_32_0_1_96_2393_out)
  );
  delay_fixed_32_0_1_1357 delay_fixed_32_0_1_1357_2394 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2412:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3203),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1357_2394_out)
  );
  delay_fixed_32_0_1_1261 delay_fixed_32_0_1_1261_2395 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2413:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3199),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1261_2395_out)
  );
  delay_fixed_32_0_1_48 delay_fixed_32_0_1_48_2396 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2414:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1340__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1486:116
    .out   (_delay_fixed_32_0_1_48_2396_out)
  );
  delay_fixed_32_0_1_1293 delay_fixed_32_0_1_1293_2397 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2415:150
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_3188),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_1293_2397_out)
  );
  delay_fixed_32_0_1_1120 delay_fixed_32_0_1_1120_2398 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2416:150
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_3184),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_1120_2398_out)
  );
  delay_fixed_32_0_1_11 delay_fixed_32_0_1_11_2399 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2417:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1330__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1476:116
    .out   (_delay_fixed_32_0_1_11_2399_out)
  );
  delay_fixed_32_0_1_1291 delay_fixed_32_0_1_1291_2400 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2418:150
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_3176),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_1291_2400_out)
  );
  delay_fixed_32_0_1_1149 delay_fixed_32_0_1_1149_2401 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2419:150
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_3172),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_1149_2401_out)
  );
  delay_fixed_32_0_1_11 delay_fixed_32_0_1_11_2402 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2420:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1330__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1476:116
    .out   (_delay_fixed_32_0_1_11_2402_out)
  );
  delay_fixed_32_0_1_288 delay_fixed_32_0_1_288_2403 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2421:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1325__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1471:116
    .out   (_delay_fixed_32_0_1_288_2403_out)
  );
  delay_fixed_32_0_1_288 delay_fixed_32_0_1_288_2404 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2422:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1325__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1471:116
    .out   (_delay_fixed_32_0_1_288_2404_out)
  );
  delay_fixed_32_0_1_169 delay_fixed_32_0_1_169_2405 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2423:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1321__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1467:116
    .out   (_delay_fixed_32_0_1_169_2405_out)
  );
  delay_fixed_32_0_1_169 delay_fixed_32_0_1_169_2406 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2424:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1321__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1467:116
    .out   (_delay_fixed_32_0_1_169_2406_out)
  );
  delay_fixed_32_0_1_39 delay_fixed_32_0_1_39_2407 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2425:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1318__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1464:116
    .out   (_delay_fixed_32_0_1_39_2407_out)
  );
  delay_fixed_32_0_1_39 delay_fixed_32_0_1_39_2408 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2426:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1318__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1464:116
    .out   (_delay_fixed_32_0_1_39_2408_out)
  );
  delay_fixed_32_0_1_11 delay_fixed_32_0_1_11_2409 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2427:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1313__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1459:116
    .out   (_delay_fixed_32_0_1_11_2409_out)
  );
  delay_fixed_32_0_1_11 delay_fixed_32_0_1_11_2410 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2428:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1313__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1459:116
    .out   (_delay_fixed_32_0_1_11_2410_out)
  );
  delay_fixed_32_0_1_175 delay_fixed_32_0_1_175_2411 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2429:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1310__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1456:136
    .out   (_delay_fixed_32_0_1_175_2411_out)
  );
  delay_fixed_32_0_1_839 delay_fixed_32_0_1_839_2412 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2430:146
    .clock (clock),
    .reset (reset),
    .in    (_dup49_const_fix_32_0_1__0000000000000235_3048),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
    .out   (_delay_fixed_32_0_1_839_2412_out)
  );
  delay_fixed_32_0_1_341 delay_fixed_32_0_1_341_2413 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2431:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1306__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1452:136
    .out   (_delay_fixed_32_0_1_341_2413_out)
  );
  delay_fixed_32_0_1_622 delay_fixed_32_0_1_622_2414 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2432:146
    .clock (clock),
    .reset (reset),
    .in    (_dup45_const_fix_32_0_1__0000000000000235_3048),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
    .out   (_delay_fixed_32_0_1_622_2414_out)
  );
  delay_fixed_32_0_1_768 delay_fixed_32_0_1_768_2415 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2433:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_3116),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_768_2415_out)
  );
  delay_fixed_32_0_1_869 delay_fixed_32_0_1_869_2416 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2434:146
    .clock (clock),
    .reset (reset),
    .in    (_dup43_const_fix_32_0_1__0000000000000235_3048),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
    .out   (_delay_fixed_32_0_1_869_2416_out)
  );
  delay_fixed_32_0_1_161 delay_fixed_32_0_1_161_2417 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2435:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1302__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1448:116
    .out   (_delay_fixed_32_0_1_161_2417_out)
  );
  delay_fixed_32_0_1_12 delay_fixed_32_0_1_12_2418 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2436:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1298__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1444:116
    .out   (_delay_fixed_32_0_1_12_2418_out)
  );
  delay_fixed_32_0_1_12 delay_fixed_32_0_1_12_2419 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2437:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1298__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1444:116
    .out   (_delay_fixed_32_0_1_12_2419_out)
  );
  delay_fixed_32_0_1_71 delay_fixed_32_0_1_71_2420 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2438:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL1294__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1440:136
    .out   (_delay_fixed_32_0_1_71_2420_out)
  );
  delay_fixed_32_0_1_719 delay_fixed_32_0_1_719_2421 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2439:146
    .clock (clock),
    .reset (reset),
    .in    (_dup33_const_fix_32_0_1__0000000000000235_3048),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
    .out   (_delay_fixed_32_0_1_719_2421_out)
  );
  delay_fixed_32_0_1_130 delay_fixed_32_0_1_130_2422 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2440:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1290__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1436:136
    .out   (_delay_fixed_32_0_1_130_2422_out)
  );
  delay_fixed_32_0_1_670 delay_fixed_32_0_1_670_2423 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2441:146
    .clock (clock),
    .reset (reset),
    .in    (_dup29_const_fix_32_0_1__0000000000000235_3048),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
    .out   (_delay_fixed_32_0_1_670_2423_out)
  );
  delay_fixed_32_0_1_678 delay_fixed_32_0_1_678_2424 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2442:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_3080),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_678_2424_out)
  );
  delay_fixed_32_0_1_781 delay_fixed_32_0_1_781_2425 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2443:146
    .clock (clock),
    .reset (reset),
    .in    (_dup27_const_fix_32_0_1__0000000000000235_3048),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
    .out   (_delay_fixed_32_0_1_781_2425_out)
  );
  delay_fixed_32_0_1_9 delay_fixed_32_0_1_9_2426 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2444:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1286__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1432:116
    .out   (_delay_fixed_32_0_1_9_2426_out)
  );
  delay_fixed_32_0_1_36 delay_fixed_32_0_1_36_2427 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2445:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL1282__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1428:136
    .out   (_delay_fixed_32_0_1_36_2427_out)
  );
  delay_fixed_32_0_1_776 delay_fixed_32_0_1_776_2428 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2446:146
    .clock (clock),
    .reset (reset),
    .in    (_dup21_const_fix_32_0_1__0000000000000235_3048),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
    .out   (_delay_fixed_32_0_1_776_2428_out)
  );
  delay_fixed_32_0_1_80 delay_fixed_32_0_1_80_2429 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2447:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL1278__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1424:136
    .out   (_delay_fixed_32_0_1_80_2429_out)
  );
  delay_fixed_32_0_1_729 delay_fixed_32_0_1_729_2430 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2448:146
    .clock (clock),
    .reset (reset),
    .in    (_dup17_const_fix_32_0_1__0000000000000235_3048),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
    .out   (_delay_fixed_32_0_1_729_2430_out)
  );
  delay_fixed_32_0_1_711 delay_fixed_32_0_1_711_2431 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2449:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_3052),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_711_2431_out)
  );
  delay_fixed_32_0_1_744 delay_fixed_32_0_1_744_2432 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2450:146
    .clock (clock),
    .reset (reset),
    .in    (_dup15_const_fix_32_0_1__0000000000000235_3048),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
    .out   (_delay_fixed_32_0_1_744_2432_out)
  );
  delay_fixed_32_0_1_3 delay_fixed_32_0_1_3_2433 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2451:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1273__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1419:116
    .out   (_delay_fixed_32_0_1_3_2433_out)
  );
  delay_fixed_32_0_1_835 delay_fixed_32_0_1_835_2434 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2452:146
    .clock (clock),
    .reset (reset),
    .in    (_dup821_const_fix_32_0_1__0000000000002000_3042),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:967:473
    .out   (_delay_fixed_32_0_1_835_2434_out)
  );
  delay_fixed_1_0_0_13 delay_fixed_1_0_0_13_2435 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2453:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1259__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1405:139
    .out   (_delay_fixed_1_0_0_13_2435_out)
  );
  delay_fixed_32_0_1_1775 delay_fixed_32_0_1_1775_2436 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2454:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2993),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1775_2436_out)
  );
  delay_fixed_32_0_1_1727 delay_fixed_32_0_1_1727_2437 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2455:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2989),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1727_2437_out)
  );
  delay_fixed_32_0_1_27 delay_fixed_32_0_1_27_2438 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2456:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1256__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1402:154
    .out   (_delay_fixed_32_0_1_27_2438_out)
  );
  delay_fixed_32_0_1_1788 delay_fixed_32_0_1_1788_2439 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2457:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2993),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1788_2439_out)
  );
  delay_fixed_32_0_1_1761 delay_fixed_32_0_1_1761_2440 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2458:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2989),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1761_2440_out)
  );
  delay_fixed_32_0_1_102 delay_fixed_32_0_1_102_2441 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2459:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1190__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1336:116
    .out   (_delay_fixed_32_0_1_102_2441_out)
  );
  delay_fixed_1_0_0_75 delay_fixed_1_0_0_75_2442 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2460:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1251__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1397:139
    .out   (_delay_fixed_1_0_0_75_2442_out)
  );
  delay_fixed_32_0_1_2017 delay_fixed_32_0_1_2017_2443 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2461:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2971),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_2017_2443_out)
  );
  delay_fixed_32_0_1_1881 delay_fixed_32_0_1_1881_2444 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2462:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2967),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1881_2444_out)
  );
  delay_fixed_32_0_1_57 delay_fixed_32_0_1_57_2445 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2463:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1248__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1394:154
    .out   (_delay_fixed_32_0_1_57_2445_out)
  );
  delay_fixed_32_0_1_1972 delay_fixed_32_0_1_1972_2446 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2464:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2971),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1972_2446_out)
  );
  delay_fixed_32_0_1_1915 delay_fixed_32_0_1_1915_2447 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2465:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2967),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1915_2447_out)
  );
  delay_fixed_32_0_1_295 delay_fixed_32_0_1_295_2448 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2466:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1200__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1346:116
    .out   (_delay_fixed_32_0_1_295_2448_out)
  );
  delay_fixed_1_0_0_20 delay_fixed_1_0_0_20_2449 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2467:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1243__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1389:139
    .out   (_delay_fixed_1_0_0_20_2449_out)
  );
  delay_fixed_32_0_1_1941 delay_fixed_32_0_1_1941_2450 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2468:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2949),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1941_2450_out)
  );
  delay_fixed_32_0_1_1846 delay_fixed_32_0_1_1846_2451 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2469:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2945),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1846_2451_out)
  );
  delay_fixed_32_0_1_50 delay_fixed_32_0_1_50_2452 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2470:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1240__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1386:154
    .out   (_delay_fixed_32_0_1_50_2452_out)
  );
  delay_fixed_32_0_1_1930 delay_fixed_32_0_1_1930_2453 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2471:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2949),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1930_2453_out)
  );
  delay_fixed_32_0_1_1880 delay_fixed_32_0_1_1880_2454 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2472:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2945),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1880_2454_out)
  );
  delay_fixed_32_0_1_356 delay_fixed_32_0_1_356_2455 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2473:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1210__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1356:116
    .out   (_delay_fixed_32_0_1_356_2455_out)
  );
  delay_fixed_1_0_0_7 delay_fixed_1_0_0_7_2456 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2474:134
    .clock (clock),
    .reset (reset),
    .in    (_LT1235__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1381:139
    .out   (_delay_fixed_1_0_0_7_2456_out)
  );
  delay_fixed_32_0_1_1774 delay_fixed_32_0_1_1774_2457 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2475:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2927),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1774_2457_out)
  );
  delay_fixed_32_0_1_1688 delay_fixed_32_0_1_1688_2458 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2476:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1688_2458_out)
  );
  delay_fixed_32_0_1_39 delay_fixed_32_0_1_39_2459 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2477:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1232__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1378:154
    .out   (_delay_fixed_32_0_1_39_2459_out)
  );
  delay_fixed_32_0_1_1761 delay_fixed_32_0_1_1761_2460 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2478:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2927),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1761_2460_out)
  );
  delay_fixed_32_0_1_1722 delay_fixed_32_0_1_1722_2461 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2479:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2923),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1722_2461_out)
  );
  delay_fixed_32_0_1_103 delay_fixed_32_0_1_103_2462 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2480:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1221__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1367:116
    .out   (_delay_fixed_32_0_1_103_2462_out)
  );
  delay_fixed_1_0_0_76 delay_fixed_1_0_0_76_2463 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2481:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1227__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1373:139
    .out   (_delay_fixed_1_0_0_76_2463_out)
  );
  delay_fixed_32_0_1_1759 delay_fixed_32_0_1_1759_2464 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2482:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2905),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1759_2464_out)
  );
  delay_fixed_32_0_1_1602 delay_fixed_32_0_1_1602_2465 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2483:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2901),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1602_2465_out)
  );
  delay_fixed_32_0_1_85 delay_fixed_32_0_1_85_2466 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2484:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1224__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1370:154
    .out   (_delay_fixed_32_0_1_85_2466_out)
  );
  delay_fixed_32_0_1_1721 delay_fixed_32_0_1_1721_2467 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2485:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2905),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1721_2467_out)
  );
  delay_fixed_32_0_1_1636 delay_fixed_32_0_1_1636_2468 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2486:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2901),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1636_2468_out)
  );
  delay_fixed_32_0_1_103 delay_fixed_32_0_1_103_2469 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2487:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1221__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1367:116
    .out   (_delay_fixed_32_0_1_103_2469_out)
  );
  delay_fixed_1_0_0_80 delay_fixed_1_0_0_80_2470 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2488:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1217__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1363:139
    .out   (_delay_fixed_1_0_0_80_2470_out)
  );
  delay_fixed_32_0_1_1918 delay_fixed_32_0_1_1918_2471 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2489:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2883),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1918_2471_out)
  );
  delay_fixed_32_0_1_1791 delay_fixed_32_0_1_1791_2472 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2490:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2879),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1791_2472_out)
  );
  delay_fixed_32_0_1_44 delay_fixed_32_0_1_44_2473 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2491:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1214__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1360:154
    .out   (_delay_fixed_32_0_1_44_2473_out)
  );
  delay_fixed_32_0_1_1869 delay_fixed_32_0_1_1869_2474 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2492:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2883),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1869_2474_out)
  );
  delay_fixed_32_0_1_1825 delay_fixed_32_0_1_1825_2475 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2493:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2879),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1825_2475_out)
  );
  delay_fixed_32_0_1_356 delay_fixed_32_0_1_356_2476 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2494:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1210__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1356:116
    .out   (_delay_fixed_32_0_1_356_2476_out)
  );
  delay_fixed_1_0_0_81 delay_fixed_1_0_0_81_2477 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2495:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1207__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1353:139
    .out   (_delay_fixed_1_0_0_81_2477_out)
  );
  delay_fixed_32_0_1_1876 delay_fixed_32_0_1_1876_2478 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2496:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2861),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1876_2478_out)
  );
  delay_fixed_32_0_1_1792 delay_fixed_32_0_1_1792_2479 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2497:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2857),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1792_2479_out)
  );
  delay_fixed_32_0_1_1 delay_fixed_32_0_1_1_2480 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2498:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1204__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1350:154
    .out   (_delay_fixed_32_0_1_1_2480_out)
  );
  delay_fixed_32_0_1_1827 delay_fixed_32_0_1_1827_2481 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2499:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2861),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1827_2481_out)
  );
  delay_fixed_32_0_1_1826 delay_fixed_32_0_1_1826_2482 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2500:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2857),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1826_2482_out)
  );
  delay_fixed_32_0_1_295 delay_fixed_32_0_1_295_2483 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2501:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1200__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1346:116
    .out   (_delay_fixed_32_0_1_295_2483_out)
  );
  delay_fixed_1_0_0_13 delay_fixed_1_0_0_13_2484 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2502:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1197__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1343:139
    .out   (_delay_fixed_1_0_0_13_2484_out)
  );
  delay_fixed_32_0_1_1798 delay_fixed_32_0_1_1798_2485 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2503:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2839),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1798_2485_out)
  );
  delay_fixed_32_0_1_1692 delay_fixed_32_0_1_1692_2486 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2504:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2835),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1692_2486_out)
  );
  delay_fixed_32_0_1_92 delay_fixed_32_0_1_92_2487 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2505:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1194__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1340:154
    .out   (_delay_fixed_32_0_1_92_2487_out)
  );
  delay_fixed_32_0_1_1818 delay_fixed_32_0_1_1818_2488 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2506:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2839),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1818_2488_out)
  );
  delay_fixed_32_0_1_1726 delay_fixed_32_0_1_1726_2489 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2507:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2835),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1726_2489_out)
  );
  delay_fixed_32_0_1_102 delay_fixed_32_0_1_102_2490 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2508:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1190__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1336:116
    .out   (_delay_fixed_32_0_1_102_2490_out)
  );
  delay_fixed_32_0_1_1679 delay_fixed_32_0_1_1679_2491 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2509:150
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_2824),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_1679_2491_out)
  );
  delay_fixed_32_0_1_1556 delay_fixed_32_0_1_1556_2492 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2510:150
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_2820),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_1556_2492_out)
  );
  delay_fixed_32_0_1_111 delay_fixed_32_0_1_111_2493 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2511:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1181__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1327:116
    .out   (_delay_fixed_32_0_1_111_2493_out)
  );
  delay_fixed_32_0_1_1687 delay_fixed_32_0_1_1687_2494 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2512:150
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_2812),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_1687_2494_out)
  );
  delay_fixed_32_0_1_1578 delay_fixed_32_0_1_1578_2495 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2513:150
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_2808),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_1578_2495_out)
  );
  delay_fixed_32_0_1_111 delay_fixed_32_0_1_111_2496 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2514:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1181__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1327:116
    .out   (_delay_fixed_32_0_1_111_2496_out)
  );
  delay_fixed_32_0_1_172 delay_fixed_32_0_1_172_2497 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2515:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1176__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1322:116
    .out   (_delay_fixed_32_0_1_172_2497_out)
  );
  delay_fixed_32_0_1_172 delay_fixed_32_0_1_172_2498 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2516:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1176__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1322:116
    .out   (_delay_fixed_32_0_1_172_2498_out)
  );
  delay_fixed_32_0_1_270 delay_fixed_32_0_1_270_2499 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2517:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1172__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1318:116
    .out   (_delay_fixed_32_0_1_270_2499_out)
  );
  delay_fixed_32_0_1_270 delay_fixed_32_0_1_270_2500 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2518:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1172__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1318:116
    .out   (_delay_fixed_32_0_1_270_2500_out)
  );
  delay_fixed_32_0_1_25 delay_fixed_32_0_1_25_2501 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2519:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1168__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1314:116
    .out   (_delay_fixed_32_0_1_25_2501_out)
  );
  delay_fixed_32_0_1_25 delay_fixed_32_0_1_25_2502 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2520:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1168__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1314:116
    .out   (_delay_fixed_32_0_1_25_2502_out)
  );
  delay_fixed_32_0_1_1 delay_fixed_32_0_1_1_2503 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2521:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1165__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1311:116
    .out   (_delay_fixed_32_0_1_1_2503_out)
  );
  delay_fixed_32_0_1_1 delay_fixed_32_0_1_1_2504 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2522:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1165__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1311:116
    .out   (_delay_fixed_32_0_1_1_2504_out)
  );
  delay_fixed_32_0_1_167 delay_fixed_32_0_1_167_2505 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2523:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1161__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1307:136
    .out   (_delay_fixed_32_0_1_167_2505_out)
  );
  delay_fixed_32_0_1_1043 delay_fixed_32_0_1_1043_2506 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2524:150
    .clock (clock),
    .reset (reset),
    .in    (_dup49_const_fix_32_0_1__0000000000000235_2684),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
    .out   (_delay_fixed_32_0_1_1043_2506_out)
  );
  delay_fixed_32_0_1_123 delay_fixed_32_0_1_123_2507 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2525:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1157__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1303:136
    .out   (_delay_fixed_32_0_1_123_2507_out)
  );
  delay_fixed_32_0_1_994 delay_fixed_32_0_1_994_2508 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2526:146
    .clock (clock),
    .reset (reset),
    .in    (_dup45_const_fix_32_0_1__0000000000000235_2684),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
    .out   (_delay_fixed_32_0_1_994_2508_out)
  );
  delay_fixed_32_0_1_986 delay_fixed_32_0_1_986_2509 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2527:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_2752),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_986_2509_out)
  );
  delay_fixed_32_0_1_1062 delay_fixed_32_0_1_1062_2510 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2528:150
    .clock (clock),
    .reset (reset),
    .in    (_dup43_const_fix_32_0_1__0000000000000235_2684),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
    .out   (_delay_fixed_32_0_1_1062_2510_out)
  );
  delay_fixed_32_0_1_7 delay_fixed_32_0_1_7_2511 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2529:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1152__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1298:116
    .out   (_delay_fixed_32_0_1_7_2511_out)
  );
  delay_fixed_32_0_1_122 delay_fixed_32_0_1_122_2512 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2530:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1149__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1295:116
    .out   (_delay_fixed_32_0_1_122_2512_out)
  );
  delay_fixed_32_0_1_920 delay_fixed_32_0_1_920_2513 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2531:146
    .clock (clock),
    .reset (reset),
    .in    (_dup29_const_fix_32_0_1__0000000000000235_2684),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
    .out   (_delay_fixed_32_0_1_920_2513_out)
  );
  delay_fixed_32_0_1_1009 delay_fixed_32_0_1_1009_2514 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2532:150
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_2716),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_1009_2514_out)
  );
  delay_fixed_32_0_1_1032 delay_fixed_32_0_1_1032_2515 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2533:150
    .clock (clock),
    .reset (reset),
    .in    (_dup27_const_fix_32_0_1__0000000000000235_2684),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
    .out   (_delay_fixed_32_0_1_1032_2515_out)
  );
  delay_fixed_32_0_1_73 delay_fixed_32_0_1_73_2516 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2534:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1137__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1283:116
    .out   (_delay_fixed_32_0_1_73_2516_out)
  );
  delay_fixed_32_0_1_138 delay_fixed_32_0_1_138_2517 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2535:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1133__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1279:136
    .out   (_delay_fixed_32_0_1_138_2517_out)
  );
  delay_fixed_32_0_1_980 delay_fixed_32_0_1_980_2518 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2536:146
    .clock (clock),
    .reset (reset),
    .in    (_dup21_const_fix_32_0_1__0000000000000235_2684),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
    .out   (_delay_fixed_32_0_1_980_2518_out)
  );
  delay_fixed_32_0_1_295 delay_fixed_32_0_1_295_2519 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2537:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1129__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1275:136
    .out   (_delay_fixed_32_0_1_295_2519_out)
  );
  delay_fixed_32_0_1_781 delay_fixed_32_0_1_781_2520 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2538:146
    .clock (clock),
    .reset (reset),
    .in    (_dup17_const_fix_32_0_1__0000000000000235_2684),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
    .out   (_delay_fixed_32_0_1_781_2520_out)
  );
  delay_fixed_32_0_1_983 delay_fixed_32_0_1_983_2521 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2539:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_2688),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_983_2521_out)
  );
  delay_fixed_32_0_1_1014 delay_fixed_32_0_1_1014_2522 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2540:150
    .clock (clock),
    .reset (reset),
    .in    (_dup15_const_fix_32_0_1__0000000000000235_2684),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
    .out   (_delay_fixed_32_0_1_1014_2522_out)
  );
  delay_fixed_32_0_1_155 delay_fixed_32_0_1_155_2523 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2541:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1124__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1270:116
    .out   (_delay_fixed_32_0_1_155_2523_out)
  );
  delay_fixed_32_0_1_915 delay_fixed_32_0_1_915_2524 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2542:146
    .clock (clock),
    .reset (reset),
    .in    (_dup821_const_fix_32_0_1__0000000000002000_2678),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:967:473
    .out   (_delay_fixed_32_0_1_915_2524_out)
  );
  delay_fixed_1_0_0_95 delay_fixed_1_0_0_95_2525 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2543:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1110__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1256:139
    .out   (_delay_fixed_1_0_0_95_2525_out)
  );
  delay_fixed_32_0_1_1777 delay_fixed_32_0_1_1777_2526 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2544:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2629),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1777_2526_out)
  );
  delay_fixed_32_0_1_1644 delay_fixed_32_0_1_1644_2527 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2545:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2625),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1644_2527_out)
  );
  delay_fixed_32_0_1_39 delay_fixed_32_0_1_39_2528 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2546:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1107__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1253:154
    .out   (_delay_fixed_32_0_1_39_2528_out)
  );
  delay_fixed_32_0_1_1717 delay_fixed_32_0_1_1717_2529 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2547:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2629),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1717_2529_out)
  );
  delay_fixed_32_0_1_1678 delay_fixed_32_0_1_1678_2530 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2548:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2625),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1678_2530_out)
  );
  delay_fixed_32_0_1_59 delay_fixed_32_0_1_59_2531 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2549:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1041__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1187:116
    .out   (_delay_fixed_32_0_1_59_2531_out)
  );
  delay_fixed_1_0_0_9 delay_fixed_1_0_0_9_2532 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2550:134
    .clock (clock),
    .reset (reset),
    .in    (_LT1102__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1248:139
    .out   (_delay_fixed_1_0_0_9_2532_out)
  );
  delay_fixed_32_0_1_2086 delay_fixed_32_0_1_2086_2533 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2551:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2607),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_2086_2533_out)
  );
  delay_fixed_32_0_1_2044 delay_fixed_32_0_1_2044_2534 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2552:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2603),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_2044_2534_out)
  );
  delay_fixed_32_0_1_7 delay_fixed_32_0_1_7_2535 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2553:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1099__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1245:154
    .out   (_delay_fixed_32_0_1_7_2535_out)
  );
  delay_fixed_32_0_1_2085 delay_fixed_32_0_1_2085_2536 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2554:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2607),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_2085_2536_out)
  );
  delay_fixed_32_0_1_2078 delay_fixed_32_0_1_2078_2537 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2555:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2603),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_2078_2537_out)
  );
  delay_fixed_32_0_1_478 delay_fixed_32_0_1_478_2538 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2556:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1051__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1197:116
    .out   (_delay_fixed_32_0_1_478_2538_out)
  );
  delay_fixed_32_0_1_2139 delay_fixed_32_0_1_2139_2539 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2557:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2493),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_2139_2539_out)
  );
  delay_fixed_32_0_1_89 delay_fixed_32_0_1_89_2540 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2558:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1055__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1201:154
    .out   (_delay_fixed_32_0_1_89_2540_out)
  );
  delay_fixed_32_0_1_2262 delay_fixed_32_0_1_2262_2541 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2559:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2497),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_2262_2541_out)
  );
  delay_fixed_32_0_1_2173 delay_fixed_32_0_1_2173_2542 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2560:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2493),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_2173_2542_out)
  );
  delay_fixed_32_0_1_478 delay_fixed_32_0_1_478_2543 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2561:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1051__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1197:116
    .out   (_delay_fixed_32_0_1_478_2543_out)
  );
  delay_fixed_1_0_0_75 delay_fixed_1_0_0_75_2544 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2562:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1048__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1194:139
    .out   (_delay_fixed_1_0_0_75_2544_out)
  );
  delay_fixed_32_0_1_1807 delay_fixed_32_0_1_1807_2545 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2563:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2475),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1807_2545_out)
  );
  delay_fixed_32_0_1_1713 delay_fixed_32_0_1_1713_2546 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2564:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2471),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1713_2546_out)
  );
  delay_fixed_32_0_1_39 delay_fixed_32_0_1_39_2547 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2565:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1045__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1191:154
    .out   (_delay_fixed_32_0_1_39_2547_out)
  );
  delay_fixed_32_0_1_1786 delay_fixed_32_0_1_1786_2548 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2566:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2475),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1786_2548_out)
  );
  delay_fixed_32_0_1_1747 delay_fixed_32_0_1_1747_2549 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2567:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2471),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1747_2549_out)
  );
  delay_fixed_32_0_1_59 delay_fixed_32_0_1_59_2550 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2568:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1041__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1187:116
    .out   (_delay_fixed_32_0_1_59_2550_out)
  );
  delay_fixed_32_0_1_1811 delay_fixed_32_0_1_1811_2551 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2569:150
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_2460),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_1811_2551_out)
  );
  delay_fixed_32_0_1_1732 delay_fixed_32_0_1_1732_2552 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2570:150
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_2456),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_1732_2552_out)
  );
  delay_fixed_32_0_1_80 delay_fixed_32_0_1_80_2553 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2571:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1032__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1178:116
    .out   (_delay_fixed_32_0_1_80_2553_out)
  );
  delay_fixed_32_0_1_1838 delay_fixed_32_0_1_1838_2554 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2572:150
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_2448),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_1838_2554_out)
  );
  delay_fixed_32_0_1_1728 delay_fixed_32_0_1_1728_2555 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2573:150
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_2444),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_1728_2555_out)
  );
  delay_fixed_32_0_1_80 delay_fixed_32_0_1_80_2556 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2574:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1032__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1178:116
    .out   (_delay_fixed_32_0_1_80_2556_out)
  );
  delay_fixed_32_0_1_226 delay_fixed_32_0_1_226_2557 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2575:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1027__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1173:116
    .out   (_delay_fixed_32_0_1_226_2557_out)
  );
  delay_fixed_32_0_1_226 delay_fixed_32_0_1_226_2558 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2576:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1027__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1173:116
    .out   (_delay_fixed_32_0_1_226_2558_out)
  );
  delay_fixed_32_0_1_256 delay_fixed_32_0_1_256_2559 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2577:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1023__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1169:116
    .out   (_delay_fixed_32_0_1_256_2559_out)
  );
  delay_fixed_32_0_1_256 delay_fixed_32_0_1_256_2560 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2578:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1023__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1169:116
    .out   (_delay_fixed_32_0_1_256_2560_out)
  );
  delay_fixed_32_0_1_23 delay_fixed_32_0_1_23_2561 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2579:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1959__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2105:154
    .out   (_delay_fixed_32_0_1_23_2561_out)
  );
  delay_fixed_32_0_1_1715 delay_fixed_32_0_1_1715_2562 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2580:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4703),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1715_2562_out)
  );
  delay_fixed_32_0_1_24 delay_fixed_32_0_1_24_2563 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2581:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1966__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2112:116
    .out   (_delay_fixed_32_0_1_24_2563_out)
  );
  delay_fixed_32_0_1_1147 delay_fixed_32_0_1_1147_2564 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2582:150
    .clock (clock),
    .reset (reset),
    .in    (_dup15_const_fix_32_0_1__0000000000000235_2320),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
    .out   (_delay_fixed_32_0_1_1147_2564_out)
  );
  delay_fixed_32_0_1_842 delay_fixed_32_0_1_842_2565 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2583:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_1988),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_842_2565_out)
  );
  delay_fixed_32_0_1_283 delay_fixed_32_0_1_283_2566 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2584:146
    .clock (clock),
    .reset (reset),
    .in    (_dup976__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1122:111
    .out   (_delay_fixed_32_0_1_283_2566_out)
  );
  delay_fixed_32_0_1_913 delay_fixed_32_0_1_913_2567 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2585:146
    .clock (clock),
    .reset (reset),
    .in    (_dup27_const_fix_32_0_1__0000000000000235_1956),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
    .out   (_delay_fixed_32_0_1_913_2567_out)
  );
  delay_fixed_32_0_1_6 delay_fixed_32_0_1_6_2568 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2586:138
    .clock (clock),
    .reset (reset),
    .in    (_MUX1971__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2117:169
    .out   (_delay_fixed_32_0_1_6_2568_out)
  );
  delay_fixed_32_0_1_1424 delay_fixed_32_0_1_1424_2569 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2587:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4725),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1424_2569_out)
  );
  delay_fixed_32_0_1_28 delay_fixed_32_0_1_28_2570 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2588:142
    .clock (clock),
    .reset (reset),
    .in    (_dup836__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:982:111
    .out   (_delay_fixed_32_0_1_28_2570_out)
  );
  delay_fixed_32_0_1_1385 delay_fixed_32_0_1_1385_2571 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2589:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4721),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1385_2571_out)
  );
  delay_fixed_32_0_1_15 delay_fixed_32_0_1_15_2572 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2590:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1969__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2115:154
    .out   (_delay_fixed_32_0_1_15_2572_out)
  );
  delay_fixed_32_0_1_1434 delay_fixed_32_0_1_1434_2573 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2591:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4725),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1434_2573_out)
  );
  delay_fixed_32_0_1_1021 delay_fixed_32_0_1_1021_2574 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2592:150
    .clock (clock),
    .reset (reset),
    .in    (_dup821_const_fix_32_0_1__0000000000002000_2314),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:967:473
    .out   (_delay_fixed_32_0_1_1021_2574_out)
  );
  delay_fixed_32_0_1_1419 delay_fixed_32_0_1_1419_2575 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2593:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4721),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1419_2575_out)
  );
  delay_fixed_32_0_1_125 delay_fixed_32_0_1_125_2576 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2594:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL833__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:979:131
    .out   (_delay_fixed_32_0_1_125_2576_out)
  );
  delay_fixed_32_0_1_692 delay_fixed_32_0_1_692_2577 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2595:146
    .clock (clock),
    .reset (reset),
    .in    (_dup21_const_fix_32_0_1__0000000000000235_1956),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
    .out   (_delay_fixed_32_0_1_692_2577_out)
  );
  delay_fixed_32_0_1_24 delay_fixed_32_0_1_24_2578 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2596:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1966__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2112:116
    .out   (_delay_fixed_32_0_1_24_2578_out)
  );
  delay_fixed_32_0_1_60 delay_fixed_32_0_1_60_2579 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2597:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL829__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:975:131
    .out   (_delay_fixed_32_0_1_60_2579_out)
  );
  delay_fixed_32_0_1_689 delay_fixed_32_0_1_689_2580 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2598:146
    .clock (clock),
    .reset (reset),
    .in    (_dup17_const_fix_32_0_1__0000000000000235_1956),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
    .out   (_delay_fixed_32_0_1_689_2580_out)
  );
  delay_fixed_32_0_1_19 delay_fixed_32_0_1_19_2581 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2599:142
    .clock (clock),
    .reset (reset),
    .in    (_MUX1961__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2107:169
    .out   (_delay_fixed_32_0_1_19_2581_out)
  );
  delay_fixed_32_0_1_1741 delay_fixed_32_0_1_1741_2582 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2600:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4703),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1741_2582_out)
  );
  delay_fixed_32_0_1_706 delay_fixed_32_0_1_706_2583 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2601:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_1960),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_706_2583_out)
  );
  delay_fixed_32_0_1_1658 delay_fixed_32_0_1_1658_2584 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2602:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4699),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1658_2584_out)
  );
  delay_fixed_32_0_1_1692 delay_fixed_32_0_1_1692_2585 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2603:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4699),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1692_2585_out)
  );
  delay_fixed_32_0_1_744 delay_fixed_32_0_1_744_2586 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2604:146
    .clock (clock),
    .reset (reset),
    .in    (_dup15_const_fix_32_0_1__0000000000000235_1956),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
    .out   (_delay_fixed_32_0_1_744_2586_out)
  );
  delay_fixed_32_0_1_13 delay_fixed_32_0_1_13_2587 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2605:142
    .clock (clock),
    .reset (reset),
    .in    (_MUX960__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1106:163
    .out   (_delay_fixed_32_0_1_13_2587_out)
  );
  delay_fixed_32_0_1_1666 delay_fixed_32_0_1_1666_2588 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2606:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2265),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1666_2588_out)
  );
  delay_fixed_32_0_1_41 delay_fixed_32_0_1_41_2589 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2607:142
    .clock (clock),
    .reset (reset),
    .in    (_dup824__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:970:111
    .out   (_delay_fixed_32_0_1_41_2589_out)
  );
  delay_fixed_32_0_1_1570 delay_fixed_32_0_1_1570_2590 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2608:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2261),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1570_2590_out)
  );
  delay_fixed_32_0_1_346 delay_fixed_32_0_1_346_2591 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2609:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1955__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2101:116
    .out   (_delay_fixed_32_0_1_346_2591_out)
  );
  delay_fixed_32_0_1_47 delay_fixed_32_0_1_47_2592 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2610:142
    .clock (clock),
    .reset (reset),
    .in    (_dup958__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1104:148
    .out   (_delay_fixed_32_0_1_47_2592_out)
  );
  delay_fixed_32_0_1_1651 delay_fixed_32_0_1_1651_2593 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2611:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2265),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1651_2593_out)
  );
  delay_fixed_32_0_1_1604 delay_fixed_32_0_1_1604_2594 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2612:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2261),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1604_2594_out)
  );
  delay_fixed_32_0_1_825 delay_fixed_32_0_1_825_2595 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2613:146
    .clock (clock),
    .reset (reset),
    .in    (_dup821_const_fix_32_0_1__0000000000002000_1950),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:967:473
    .out   (_delay_fixed_32_0_1_825_2595_out)
  );
  delay_fixed_32_0_1_62 delay_fixed_32_0_1_62_2596 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2614:142
    .clock (clock),
    .reset (reset),
    .in    (_MUX1951__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2097:169
    .out   (_delay_fixed_32_0_1_62_2596_out)
  );
  delay_fixed_32_0_1_1702 delay_fixed_32_0_1_1702_2597 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2615:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4681),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1702_2597_out)
  );
  delay_fixed_32_0_1_190 delay_fixed_32_0_1_190_2598 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2616:146
    .clock (clock),
    .reset (reset),
    .in    (_dup890__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1036:111
    .out   (_delay_fixed_32_0_1_190_2598_out)
  );
  delay_fixed_32_0_1_1609 delay_fixed_32_0_1_1609_2599 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2617:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4677),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1609_2599_out)
  );
  delay_fixed_32_0_1_29 delay_fixed_32_0_1_29_2600 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2618:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1949__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2095:154
    .out   (_delay_fixed_32_0_1_29_2600_out)
  );
  delay_fixed_32_0_1_1672 delay_fixed_32_0_1_1672_2601 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2619:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4681),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1672_2601_out)
  );
  delay_fixed_1_0_0_53 delay_fixed_1_0_0_53_2602 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2620:138
    .clock (clock),
    .reset (reset),
    .in    (_LT953__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1099:134
    .out   (_delay_fixed_1_0_0_53_2602_out)
  );
  delay_fixed_32_0_1_1963 delay_fixed_32_0_1_1963_2603 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2621:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2243),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1963_2603_out)
  );
  delay_fixed_32_0_1_1643 delay_fixed_32_0_1_1643_2604 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2622:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4677),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1643_2604_out)
  );
  delay_fixed_32_0_1_1881 delay_fixed_32_0_1_1881_2605 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2623:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2239),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1881_2605_out)
  );
  delay_fixed_32_0_1_41 delay_fixed_32_0_1_41_2606 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2624:142
    .clock (clock),
    .reset (reset),
    .in    (_dup950__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1096:148
    .out   (_delay_fixed_32_0_1_41_2606_out)
  );
  delay_fixed_32_0_1_1956 delay_fixed_32_0_1_1956_2607 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2625:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2243),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1956_2607_out)
  );
  delay_fixed_32_0_1_1915 delay_fixed_32_0_1_1915_2608 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2626:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2239),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1915_2608_out)
  );
  delay_fixed_32_0_1_342 delay_fixed_32_0_1_342_2609 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2627:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1945__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2091:116
    .out   (_delay_fixed_32_0_1_342_2609_out)
  );
  delay_fixed_32_0_1_460 delay_fixed_32_0_1_460_2610 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2628:146
    .clock (clock),
    .reset (reset),
    .in    (_dup902__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1048:111
    .out   (_delay_fixed_32_0_1_460_2610_out)
  );
  delay_fixed_1_0_0_52 delay_fixed_1_0_0_52_2611 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2629:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1942__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2088:139
    .out   (_delay_fixed_1_0_0_52_2611_out)
  );
  delay_fixed_32_0_1_1575 delay_fixed_32_0_1_1575_2612 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2630:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4659),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1575_2612_out)
  );
  delay_fixed_32_0_1_33 delay_fixed_32_0_1_33_2613 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2631:142
    .clock (clock),
    .reset (reset),
    .in    (_MUX944__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1090:163
    .out   (_delay_fixed_32_0_1_33_2613_out)
  );
  delay_fixed_32_0_1_1758 delay_fixed_32_0_1_1758_2614 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2632:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2221),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1758_2614_out)
  );
  delay_fixed_32_0_1_1454 delay_fixed_32_0_1_1454_2615 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2633:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4655),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1454_2615_out)
  );
  delay_fixed_32_0_1_1702 delay_fixed_32_0_1_1702_2616 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2634:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2217),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1702_2616_out)
  );
  delay_fixed_32_0_1_85 delay_fixed_32_0_1_85_2617 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2635:142
    .clock (clock),
    .reset (reset),
    .in    (_dup779__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:925:111
    .out   (_delay_fixed_32_0_1_85_2617_out)
  );
  delay_fixed_32_0_1_40 delay_fixed_32_0_1_40_2618 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2636:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1939__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2085:154
    .out   (_delay_fixed_32_0_1_40_2618_out)
  );
  delay_fixed_32_0_1_1528 delay_fixed_32_0_1_1528_2619 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2637:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4659),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1528_2619_out)
  );
  delay_fixed_32_0_1_22 delay_fixed_32_0_1_22_2620 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2638:142
    .clock (clock),
    .reset (reset),
    .in    (_dup942__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1088:148
    .out   (_delay_fixed_32_0_1_22_2620_out)
  );
  delay_fixed_32_0_1_1758 delay_fixed_32_0_1_1758_2621 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2639:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2221),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1758_2621_out)
  );
  delay_fixed_32_0_1_1488 delay_fixed_32_0_1_1488_2622 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2640:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4655),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1488_2622_out)
  );
  delay_fixed_32_0_1_1736 delay_fixed_32_0_1_1736_2623 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2641:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2217),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1736_2623_out)
  );
  delay_fixed_32_0_1_149 delay_fixed_32_0_1_149_2624 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2642:146
    .clock (clock),
    .reset (reset),
    .in    (_dup784__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:930:111
    .out   (_delay_fixed_32_0_1_149_2624_out)
  );
  delay_fixed_32_0_1_39 delay_fixed_32_0_1_39_2625 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2643:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1936__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2082:116
    .out   (_delay_fixed_32_0_1_39_2625_out)
  );
  delay_fixed_32_0_1_342 delay_fixed_32_0_1_342_2626 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2644:146
    .clock (clock),
    .reset (reset),
    .in    (_dup912__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1058:111
    .out   (_delay_fixed_32_0_1_342_2626_out)
  );
  delay_fixed_32_0_1_151 delay_fixed_32_0_1_151_2627 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2645:146
    .clock (clock),
    .reset (reset),
    .in    (_dup789__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:935:111
    .out   (_delay_fixed_32_0_1_151_2627_out)
  );
  delay_fixed_32_0_1_11 delay_fixed_32_0_1_11_2628 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2646:142
    .clock (clock),
    .reset (reset),
    .in    (_MUX936__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1082:163
    .out   (_delay_fixed_32_0_1_11_2628_out)
  );
  delay_fixed_32_0_1_1575 delay_fixed_32_0_1_1575_2629 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2647:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2199),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1575_2629_out)
  );
  delay_fixed_32_0_1_1511 delay_fixed_32_0_1_1511_2630 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2648:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2195),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1511_2630_out)
  );
  delay_fixed_32_0_1_1379 delay_fixed_32_0_1_1379_2631 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2649:150
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_4644),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_1379_2631_out)
  );
  delay_fixed_32_0_1_22 delay_fixed_32_0_1_22_2632 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2650:142
    .clock (clock),
    .reset (reset),
    .in    (_dup795__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:941:111
    .out   (_delay_fixed_32_0_1_22_2632_out)
  );
  delay_fixed_32_0_1_1277 delay_fixed_32_0_1_1277_2633 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2651:150
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_4640),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_1277_2633_out)
  );
  delay_fixed_32_0_1_24 delay_fixed_32_0_1_24_2634 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2652:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1926__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2072:116
    .out   (_delay_fixed_32_0_1_24_2634_out)
  );
  delay_fixed_32_0_1_22 delay_fixed_32_0_1_22_2635 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2653:142
    .clock (clock),
    .reset (reset),
    .in    (_dup795__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:941:111
    .out   (_delay_fixed_32_0_1_22_2635_out)
  );
  delay_fixed_32_0_1_1362 delay_fixed_32_0_1_1362_2636 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2654:150
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_4632),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_1362_2636_out)
  );
  delay_fixed_32_0_1_1238 delay_fixed_32_0_1_1238_2637 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2655:150
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_4628),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_1238_2637_out)
  );
  delay_fixed_32_0_1_24 delay_fixed_32_0_1_24_2638 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2656:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1926__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2072:116
    .out   (_delay_fixed_32_0_1_24_2638_out)
  );
  delay_fixed_32_0_1_151 delay_fixed_32_0_1_151_2639 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2657:146
    .clock (clock),
    .reset (reset),
    .in    (_dup789__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:935:111
    .out   (_delay_fixed_32_0_1_151_2639_out)
  );
  delay_fixed_32_0_1_121 delay_fixed_32_0_1_121_2640 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2658:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1921__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2067:116
    .out   (_delay_fixed_32_0_1_121_2640_out)
  );
  delay_fixed_32_0_1_121 delay_fixed_32_0_1_121_2641 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2659:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1921__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2067:116
    .out   (_delay_fixed_32_0_1_121_2641_out)
  );
  delay_fixed_32_0_1_235 delay_fixed_32_0_1_235_2642 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2660:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1917__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2063:116
    .out   (_delay_fixed_32_0_1_235_2642_out)
  );
  delay_fixed_32_0_1_149 delay_fixed_32_0_1_149_2643 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2661:146
    .clock (clock),
    .reset (reset),
    .in    (_dup784__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:930:111
    .out   (_delay_fixed_32_0_1_149_2643_out)
  );
  delay_fixed_32_0_1_235 delay_fixed_32_0_1_235_2644 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2662:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1917__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2063:116
    .out   (_delay_fixed_32_0_1_235_2644_out)
  );
  delay_fixed_32_0_1_75 delay_fixed_32_0_1_75_2645 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2663:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1913__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2059:116
    .out   (_delay_fixed_32_0_1_75_2645_out)
  );
  delay_fixed_32_0_1_75 delay_fixed_32_0_1_75_2646 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2664:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1913__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2059:116
    .out   (_delay_fixed_32_0_1_75_2646_out)
  );
  delay_fixed_32_0_1_26 delay_fixed_32_0_1_26_2647 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2665:142
    .clock (clock),
    .reset (reset),
    .in    (_dup934__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1080:148
    .out   (_delay_fixed_32_0_1_26_2647_out)
  );
  delay_fixed_32_0_1_1571 delay_fixed_32_0_1_1571_2648 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2666:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2199),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1571_2648_out)
  );
  delay_fixed_32_0_1_85 delay_fixed_32_0_1_85_2649 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2667:142
    .clock (clock),
    .reset (reset),
    .in    (_dup779__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:925:111
    .out   (_delay_fixed_32_0_1_85_2649_out)
  );
  delay_fixed_32_0_1_1545 delay_fixed_32_0_1_1545_2650 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2668:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2195),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1545_2650_out)
  );
  delay_fixed_32_0_1_3 delay_fixed_32_0_1_3_2651 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2669:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1909__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2055:116
    .out   (_delay_fixed_32_0_1_3_2651_out)
  );
  delay_fixed_32_0_1_3 delay_fixed_32_0_1_3_2652 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2670:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1909__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2055:116
    .out   (_delay_fixed_32_0_1_3_2652_out)
  );
  delay_fixed_32_0_1_127 delay_fixed_32_0_1_127_2653 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2671:146
    .clock (clock),
    .reset (reset),
    .in    (_dup922__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1068:111
    .out   (_delay_fixed_32_0_1_127_2653_out)
  );
  delay_fixed_32_0_1_622 delay_fixed_32_0_1_622_2654 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2672:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_1844),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_622_2654_out)
  );
  delay_fixed_32_0_1_473 delay_fixed_32_0_1_473_2655 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2673:146
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_1840),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_473_2655_out)
  );
  delay_fixed_1_0_0_108 delay_fixed_1_0_0_108_2656 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2674:142
    .clock (clock),
    .reset (reset),
    .in    (_LT929__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1075:134
    .out   (_delay_fixed_1_0_0_108_2656_out)
  );
  delay_fixed_32_0_1_1550 delay_fixed_32_0_1_1550_2657 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2675:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2177),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1550_2657_out)
  );
  delay_fixed_32_0_1_12 delay_fixed_32_0_1_12_2658 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2676:142
    .clock (clock),
    .reset (reset),
    .in    (_dup769__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:915:111
    .out   (_delay_fixed_32_0_1_12_2658_out)
  );
  delay_fixed_32_0_1_1399 delay_fixed_32_0_1_1399_2659 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2677:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2173),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1399_2659_out)
  );
  delay_fixed_32_0_1_174 delay_fixed_32_0_1_174_2660 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2678:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1906__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2052:136
    .out   (_delay_fixed_32_0_1_174_2660_out)
  );
  delay_fixed_32_0_1_96 delay_fixed_32_0_1_96_2661 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2679:142
    .clock (clock),
    .reset (reset),
    .in    (_dup926__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1072:148
    .out   (_delay_fixed_32_0_1_96_2661_out)
  );
  delay_fixed_32_0_1_1529 delay_fixed_32_0_1_1529_2662 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2680:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2177),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1529_2662_out)
  );
  delay_fixed_32_0_1_552 delay_fixed_32_0_1_552_2663 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2681:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_1832),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_552_2663_out)
  );
  delay_fixed_32_0_1_732 delay_fixed_32_0_1_732_2664 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2682:146
    .clock (clock),
    .reset (reset),
    .in    (_dup49_const_fix_32_0_1__0000000000000235_4504),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
    .out   (_delay_fixed_32_0_1_732_2664_out)
  );
  delay_fixed_32_0_1_1433 delay_fixed_32_0_1_1433_2665 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2683:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2173),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1433_2665_out)
  );
  delay_fixed_32_0_1_472 delay_fixed_32_0_1_472_2666 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2684:146
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_1828),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_472_2666_out)
  );
  delay_fixed_32_0_1_12 delay_fixed_32_0_1_12_2667 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2685:142
    .clock (clock),
    .reset (reset),
    .in    (_dup769__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:915:111
    .out   (_delay_fixed_32_0_1_12_2667_out)
  );
  delay_fixed_32_0_1_195 delay_fixed_32_0_1_195_2668 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2686:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1902__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2048:136
    .out   (_delay_fixed_32_0_1_195_2668_out)
  );
  delay_fixed_32_0_1_127 delay_fixed_32_0_1_127_2669 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2687:146
    .clock (clock),
    .reset (reset),
    .in    (_dup922__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1068:111
    .out   (_delay_fixed_32_0_1_127_2669_out)
  );
  delay_fixed_32_0_1_673 delay_fixed_32_0_1_673_2670 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2688:146
    .clock (clock),
    .reset (reset),
    .in    (_dup45_const_fix_32_0_1__0000000000000235_4504),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
    .out   (_delay_fixed_32_0_1_673_2670_out)
  );
  delay_fixed_32_0_1_50 delay_fixed_32_0_1_50_2671 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2689:142
    .clock (clock),
    .reset (reset),
    .in    (_dup765__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:911:111
    .out   (_delay_fixed_32_0_1_50_2671_out)
  );
  delay_fixed_32_0_1_658 delay_fixed_32_0_1_658_2672 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2690:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_4572),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_658_2672_out)
  );
  delay_fixed_32_0_1_50 delay_fixed_32_0_1_50_2673 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2691:142
    .clock (clock),
    .reset (reset),
    .in    (_dup765__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:911:111
    .out   (_delay_fixed_32_0_1_50_2673_out)
  );
  delay_fixed_32_0_1_769 delay_fixed_32_0_1_769_2674 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2692:146
    .clock (clock),
    .reset (reset),
    .in    (_dup43_const_fix_32_0_1__0000000000000235_4504),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
    .out   (_delay_fixed_32_0_1_769_2674_out)
  );
  delay_fixed_32_0_1_3 delay_fixed_32_0_1_3_2675 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2693:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1898__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2044:116
    .out   (_delay_fixed_32_0_1_3_2675_out)
  );
  delay_fixed_1_0_0_27 delay_fixed_1_0_0_27_2676 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2694:138
    .clock (clock),
    .reset (reset),
    .in    (_LT919__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1065:134
    .out   (_delay_fixed_1_0_0_27_2676_out)
  );
  delay_fixed_32_0_1_1781 delay_fixed_32_0_1_1781_2677 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2695:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2155),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1781_2677_out)
  );
  delay_fixed_32_0_1_1716 delay_fixed_32_0_1_1716_2678 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2696:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2151),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1716_2678_out)
  );
  delay_fixed_32_0_1_55 delay_fixed_32_0_1_55_2679 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2697:142
    .clock (clock),
    .reset (reset),
    .in    (_dup761__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:907:111
    .out   (_delay_fixed_32_0_1_55_2679_out)
  );
  delay_fixed_32_0_1_19 delay_fixed_32_0_1_19_2680 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2698:142
    .clock (clock),
    .reset (reset),
    .in    (_dup916__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1062:148
    .out   (_delay_fixed_32_0_1_19_2680_out)
  );
  delay_fixed_32_0_1_1769 delay_fixed_32_0_1_1769_2681 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2699:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2155),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1769_2681_out)
  );
  delay_fixed_32_0_1_55 delay_fixed_32_0_1_55_2682 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2700:142
    .clock (clock),
    .reset (reset),
    .in    (_dup761__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:907:111
    .out   (_delay_fixed_32_0_1_55_2682_out)
  );
  delay_fixed_32_0_1_29 delay_fixed_32_0_1_29_2683 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2701:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1893__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2039:116
    .out   (_delay_fixed_32_0_1_29_2683_out)
  );
  delay_fixed_32_0_1_1750 delay_fixed_32_0_1_1750_2684 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2702:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2151),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1750_2684_out)
  );
  delay_fixed_32_0_1_29 delay_fixed_32_0_1_29_2685 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2703:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1893__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2039:116
    .out   (_delay_fixed_32_0_1_29_2685_out)
  );
  delay_fixed_32_0_1_1 delay_fixed_32_0_1_1_2686 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2704:138
    .clock (clock),
    .reset (reset),
    .in    (_dup757__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:903:111
    .out   (_delay_fixed_32_0_1_1_2686_out)
  );
  delay_fixed_32_0_1_342 delay_fixed_32_0_1_342_2687 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2705:146
    .clock (clock),
    .reset (reset),
    .in    (_dup912__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1058:111
    .out   (_delay_fixed_32_0_1_342_2687_out)
  );
  delay_fixed_32_0_1_1 delay_fixed_32_0_1_1_2688 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2706:138
    .clock (clock),
    .reset (reset),
    .in    (_dup757__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:903:111
    .out   (_delay_fixed_32_0_1_1_2688_out)
  );
  delay_fixed_32_0_1_313 delay_fixed_32_0_1_313_2689 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2707:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1890__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2036:136
    .out   (_delay_fixed_32_0_1_313_2689_out)
  );
  delay_fixed_32_0_1_652 delay_fixed_32_0_1_652_2690 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2708:146
    .clock (clock),
    .reset (reset),
    .in    (_dup33_const_fix_32_0_1__0000000000000235_4504),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
    .out   (_delay_fixed_32_0_1_652_2690_out)
  );
  delay_fixed_32_0_1_135 delay_fixed_32_0_1_135_2691 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2709:146
    .clock (clock),
    .reset (reset),
    .in    (_dup754__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:900:111
    .out   (_delay_fixed_32_0_1_135_2691_out)
  );
  delay_fixed_1_0_0_36 delay_fixed_1_0_0_36_2692 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2710:138
    .clock (clock),
    .reset (reset),
    .in    (_LT909__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1055:134
    .out   (_delay_fixed_1_0_0_36_2692_out)
  );
  delay_fixed_32_0_1_1824 delay_fixed_32_0_1_1824_2693 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2711:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2133),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1824_2693_out)
  );
  delay_fixed_32_0_1_135 delay_fixed_32_0_1_135_2694 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2712:146
    .clock (clock),
    .reset (reset),
    .in    (_dup754__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:900:111
    .out   (_delay_fixed_32_0_1_135_2694_out)
  );
  delay_fixed_32_0_1_176 delay_fixed_32_0_1_176_2695 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2713:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1886__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2032:136
    .out   (_delay_fixed_32_0_1_176_2695_out)
  );
  delay_fixed_32_0_1_1726 delay_fixed_32_0_1_1726_2696 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2714:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2129),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1726_2696_out)
  );
  delay_fixed_32_0_1_27 delay_fixed_32_0_1_27_2697 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2715:142
    .clock (clock),
    .reset (reset),
    .in    (_dup906__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1052:148
    .out   (_delay_fixed_32_0_1_27_2697_out)
  );
  delay_fixed_32_0_1_1787 delay_fixed_32_0_1_1787_2698 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2716:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2133),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1787_2698_out)
  );
  delay_fixed_32_0_1_725 delay_fixed_32_0_1_725_2699 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2717:146
    .clock (clock),
    .reset (reset),
    .in    (_dup29_const_fix_32_0_1__0000000000000235_4504),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
    .out   (_delay_fixed_32_0_1_725_2699_out)
  );
  delay_fixed_32_0_1_1760 delay_fixed_32_0_1_1760_2700 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2718:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2129),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1760_2700_out)
  );
  delay_fixed_32_0_1_198 delay_fixed_32_0_1_198_2701 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2719:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL751__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:897:131
    .out   (_delay_fixed_32_0_1_198_2701_out)
  );
  delay_fixed_32_0_1_742 delay_fixed_32_0_1_742_2702 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2720:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_4536),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_742_2702_out)
  );
  delay_fixed_32_0_1_74 delay_fixed_32_0_1_74_2703 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2721:142
    .clock (clock),
    .reset (reset),
    .in    (_dup49_const_fix_32_0_1__0000000000000235_1725),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
    .out   (_delay_fixed_32_0_1_74_2703_out)
  );
  delay_fixed_32_0_1_808 delay_fixed_32_0_1_808_2704 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2722:146
    .clock (clock),
    .reset (reset),
    .in    (_dup27_const_fix_32_0_1__0000000000000235_4504),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
    .out   (_delay_fixed_32_0_1_808_2704_out)
  );
  delay_fixed_32_0_1_141 delay_fixed_32_0_1_141_2705 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2723:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL748__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:894:131
    .out   (_delay_fixed_32_0_1_141_2705_out)
  );
  delay_fixed_32_0_1_131 delay_fixed_32_0_1_131_2706 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2724:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1882__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2028:116
    .out   (_delay_fixed_32_0_1_131_2706_out)
  );
  delay_fixed_32_0_1_460 delay_fixed_32_0_1_460_2707 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2725:146
    .clock (clock),
    .reset (reset),
    .in    (_dup902__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1048:111
    .out   (_delay_fixed_32_0_1_460_2707_out)
  );
  delay_fixed_32_0_1_98 delay_fixed_32_0_1_98_2708 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2726:142
    .clock (clock),
    .reset (reset),
    .in    (_dup45_const_fix_32_0_1__0000000000000235_1725),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
    .out   (_delay_fixed_32_0_1_98_2708_out)
  );
  delay_fixed_32_0_1_155 delay_fixed_32_0_1_155_2709 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2727:146
    .clock (clock),
    .reset (reset),
    .in    (_dup43_const_fix_32_0_1__0000000000000235_1725),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
    .out   (_delay_fixed_32_0_1_155_2709_out)
  );
  delay_fixed_32_0_1_80 delay_fixed_32_0_1_80_2710 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2728:142
    .clock (clock),
    .reset (reset),
    .in    (_dup744__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:890:111
    .out   (_delay_fixed_32_0_1_80_2710_out)
  );
  delay_fixed_32_0_1_119 delay_fixed_32_0_1_119_2711 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2729:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1878__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2024:136
    .out   (_delay_fixed_32_0_1_119_2711_out)
  );
  delay_fixed_32_0_1_53 delay_fixed_32_0_1_53_2712 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2730:142
    .clock (clock),
    .reset (reset),
    .in    (_MUX897__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1043:163
    .out   (_delay_fixed_32_0_1_53_2712_out)
  );
  delay_fixed_32_0_1_1623 delay_fixed_32_0_1_1623_2713 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2731:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2111),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1623_2713_out)
  );
  delay_fixed_32_0_1_779 delay_fixed_32_0_1_779_2714 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2732:146
    .clock (clock),
    .reset (reset),
    .in    (_dup21_const_fix_32_0_1__0000000000000235_4504),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
    .out   (_delay_fixed_32_0_1_779_2714_out)
  );
  delay_fixed_32_0_1_1526 delay_fixed_32_0_1_1526_2715 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2733:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1526_2715_out)
  );
  delay_fixed_32_0_1_3 delay_fixed_32_0_1_3_2716 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2734:138
    .clock (clock),
    .reset (reset),
    .in    (_dup741__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:887:111
    .out   (_delay_fixed_32_0_1_3_2716_out)
  );
  delay_fixed_32_0_1_243 delay_fixed_32_0_1_243_2717 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2735:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1874__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2020:136
    .out   (_delay_fixed_32_0_1_243_2717_out)
  );
  delay_fixed_32_0_1_40 delay_fixed_32_0_1_40_2718 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2736:142
    .clock (clock),
    .reset (reset),
    .in    (_dup894__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1040:148
    .out   (_delay_fixed_32_0_1_40_2718_out)
  );
  delay_fixed_32_0_1_1600 delay_fixed_32_0_1_1600_2719 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2737:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2111),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1600_2719_out)
  );
  delay_fixed_32_0_1_3 delay_fixed_32_0_1_3_2720 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2738:138
    .clock (clock),
    .reset (reset),
    .in    (_dup741__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:887:111
    .out   (_delay_fixed_32_0_1_3_2720_out)
  );
  delay_fixed_32_0_1_1560 delay_fixed_32_0_1_1560_2721 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2739:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1560_2721_out)
  );
  delay_fixed_32_0_1_647 delay_fixed_32_0_1_647_2722 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2740:146
    .clock (clock),
    .reset (reset),
    .in    (_dup17_const_fix_32_0_1__0000000000000235_4504),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
    .out   (_delay_fixed_32_0_1_647_2722_out)
  );
  delay_fixed_32_0_1_805 delay_fixed_32_0_1_805_2723 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2741:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_4508),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_805_2723_out)
  );
  delay_fixed_32_0_1_17 delay_fixed_32_0_1_17_2724 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2742:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL738__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:884:131
    .out   (_delay_fixed_32_0_1_17_2724_out)
  );
  delay_fixed_32_0_1_813 delay_fixed_32_0_1_813_2725 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2743:146
    .clock (clock),
    .reset (reset),
    .in    (_dup15_const_fix_32_0_1__0000000000000235_4504),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
    .out   (_delay_fixed_32_0_1_813_2725_out)
  );
  delay_fixed_32_0_1_119 delay_fixed_32_0_1_119_2726 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2744:146
    .clock (clock),
    .reset (reset),
    .in    (_dup33_const_fix_32_0_1__0000000000000235_1725),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
    .out   (_delay_fixed_32_0_1_119_2726_out)
  );
  delay_fixed_32_0_1_88 delay_fixed_32_0_1_88_2727 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2745:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1869__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2015:116
    .out   (_delay_fixed_32_0_1_88_2727_out)
  );
  delay_fixed_32_0_1_131 delay_fixed_32_0_1_131_2728 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2746:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL735__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:881:131
    .out   (_delay_fixed_32_0_1_131_2728_out)
  );
  delay_fixed_32_0_1_21 delay_fixed_32_0_1_21_2729 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2747:142
    .clock (clock),
    .reset (reset),
    .in    (_dup731__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:877:111
    .out   (_delay_fixed_32_0_1_21_2729_out)
  );
  delay_fixed_32_0_1_765 delay_fixed_32_0_1_765_2730 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2748:146
    .clock (clock),
    .reset (reset),
    .in    (_dup821_const_fix_32_0_1__0000000000002000_4498),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:967:473
    .out   (_delay_fixed_32_0_1_765_2730_out)
  );
  delay_fixed_32_0_1_124 delay_fixed_32_0_1_124_2731 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2749:146
    .clock (clock),
    .reset (reset),
    .in    (_dup27_const_fix_32_0_1__0000000000000235_1725),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
    .out   (_delay_fixed_32_0_1_124_2731_out)
  );
  delay_fixed_32_0_1_82 delay_fixed_32_0_1_82_2732 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2750:142
    .clock (clock),
    .reset (reset),
    .in    (_dup731__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:877:111
    .out   (_delay_fixed_32_0_1_82_2732_out)
  );
  delay_fixed_32_0_1_122 delay_fixed_32_0_1_122_2733 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2751:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL729__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:875:131
    .out   (_delay_fixed_32_0_1_122_2733_out)
  );
  delay_fixed_32_0_1_53 delay_fixed_32_0_1_53_2734 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2752:142
    .clock (clock),
    .reset (reset),
    .in    (_dup21_const_fix_32_0_1__0000000000000235_1725),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
    .out   (_delay_fixed_32_0_1_53_2734_out)
  );
  delay_fixed_32_0_1_88 delay_fixed_32_0_1_88_2735 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2753:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL726__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:872:131
    .out   (_delay_fixed_32_0_1_88_2735_out)
  );
  delay_fixed_32_0_1_4 delay_fixed_32_0_1_4_2736 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2754:138
    .clock (clock),
    .reset (reset),
    .in    (_dup722__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:868:111
    .out   (_delay_fixed_32_0_1_4_2736_out)
  );
  delay_fixed_32_0_1_75 delay_fixed_32_0_1_75_2737 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2755:142
    .clock (clock),
    .reset (reset),
    .in    (_dup15_const_fix_32_0_1__0000000000000235_1725),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
    .out   (_delay_fixed_32_0_1_75_2737_out)
  );
  delay_fixed_32_0_1_13 delay_fixed_32_0_1_13_2738 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2756:142
    .clock (clock),
    .reset (reset),
    .in    (_dup722__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:868:111
    .out   (_delay_fixed_32_0_1_13_2738_out)
  );
  delay_fixed_1_0_0_32 delay_fixed_1_0_0_32_2739 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2757:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1855__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2001:139
    .out   (_delay_fixed_1_0_0_32_2739_out)
  );
  delay_fixed_32_0_1_1597 delay_fixed_32_0_1_1597_2740 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2758:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4449),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1597_2740_out)
  );
  delay_fixed_32_0_1_1549 delay_fixed_32_0_1_1549_2741 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2759:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4445),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1549_2741_out)
  );
  delay_fixed_32_0_1_134 delay_fixed_32_0_1_134_2742 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2760:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_1719),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_134_2742_out)
  );
  delay_fixed_32_0_1_41 delay_fixed_32_0_1_41_2743 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2761:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1852__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1998:154
    .out   (_delay_fixed_32_0_1_41_2743_out)
  );
  delay_fixed_32_0_1_1624 delay_fixed_32_0_1_1624_2744 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2762:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4449),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1624_2744_out)
  );
  delay_fixed_32_0_1_1583 delay_fixed_32_0_1_1583_2745 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2763:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4445),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1583_2745_out)
  );
  delay_fixed_32_0_1_158 delay_fixed_32_0_1_158_2746 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2764:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1786__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1932:116
    .out   (_delay_fixed_32_0_1_158_2746_out)
  );
  delay_fixed_1_0_0_8 delay_fixed_1_0_0_8_2747 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2765:134
    .clock (clock),
    .reset (reset),
    .in    (_LT1847__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1993:139
    .out   (_delay_fixed_1_0_0_8_2747_out)
  );
  delay_fixed_32_0_1_1899 delay_fixed_32_0_1_1899_2748 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2766:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4427),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1899_2748_out)
  );
  delay_fixed_32_0_1_1813 delay_fixed_32_0_1_1813_2749 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2767:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4423),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1813_2749_out)
  );
  delay_fixed_32_0_1_35 delay_fixed_32_0_1_35_2750 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2768:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1844__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1990:154
    .out   (_delay_fixed_32_0_1_35_2750_out)
  );
  delay_fixed_32_0_1_1882 delay_fixed_32_0_1_1882_2751 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2769:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4427),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1882_2751_out)
  );
  delay_fixed_32_0_1_1847 delay_fixed_32_0_1_1847_2752 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2770:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4423),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1847_2752_out)
  );
  delay_fixed_32_0_1_440 delay_fixed_32_0_1_440_2753 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2771:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1796__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1942:116
    .out   (_delay_fixed_32_0_1_440_2753_out)
  );
  delay_fixed_32_0_1_90 delay_fixed_32_0_1_90_2754 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2772:142
    .clock (clock),
    .reset (reset),
    .in    (_dup680__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:826:111
    .out   (_delay_fixed_32_0_1_90_2754_out)
  );
  delay_fixed_1_0_0_60 delay_fixed_1_0_0_60_2755 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2773:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1839__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1985:139
    .out   (_delay_fixed_1_0_0_60_2755_out)
  );
  delay_fixed_32_0_1_1980 delay_fixed_32_0_1_1980_2756 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2774:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4405),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1980_2756_out)
  );
  delay_fixed_32_0_1_1902 delay_fixed_32_0_1_1902_2757 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2775:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4401),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1902_2757_out)
  );
  delay_fixed_32_0_1_65 delay_fixed_32_0_1_65_2758 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2776:142
    .clock (clock),
    .reset (reset),
    .in    (_dup684__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:830:111
    .out   (_delay_fixed_32_0_1_65_2758_out)
  );
  delay_fixed_32_0_1_32 delay_fixed_32_0_1_32_2759 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2777:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1836__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1982:154
    .out   (_delay_fixed_32_0_1_32_2759_out)
  );
  delay_fixed_32_0_1_1968 delay_fixed_32_0_1_1968_2760 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2778:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4405),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1968_2760_out)
  );
  delay_fixed_32_0_1_1936 delay_fixed_32_0_1_1936_2761 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2779:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4401),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1936_2761_out)
  );
  delay_fixed_32_0_1_249 delay_fixed_32_0_1_249_2762 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2780:146
    .clock (clock),
    .reset (reset),
    .in    (_dup689__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:835:111
    .out   (_delay_fixed_32_0_1_249_2762_out)
  );
  delay_fixed_32_0_1_445 delay_fixed_32_0_1_445_2763 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2781:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1806__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1952:116
    .out   (_delay_fixed_32_0_1_445_2763_out)
  );
  delay_fixed_32_0_1_108 delay_fixed_32_0_1_108_2764 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2782:146
    .clock (clock),
    .reset (reset),
    .in    (_dup695__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:841:111
    .out   (_delay_fixed_32_0_1_108_2764_out)
  );
  delay_fixed_1_0_0_97 delay_fixed_1_0_0_97_2765 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2783:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1831__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1977:139
    .out   (_delay_fixed_1_0_0_97_2765_out)
  );
  delay_fixed_32_0_1_1806 delay_fixed_32_0_1_1806_2766 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2784:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4383),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1806_2766_out)
  );
  delay_fixed_32_0_1_1693 delay_fixed_32_0_1_1693_2767 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2785:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4379),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1693_2767_out)
  );
  delay_fixed_32_0_1_54 delay_fixed_32_0_1_54_2768 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2786:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1828__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1974:154
    .out   (_delay_fixed_32_0_1_54_2768_out)
  );
  delay_fixed_32_0_1_1781 delay_fixed_32_0_1_1781_2769 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2787:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4383),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1781_2769_out)
  );
  delay_fixed_32_0_1_108 delay_fixed_32_0_1_108_2770 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2788:146
    .clock (clock),
    .reset (reset),
    .in    (_dup695__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:841:111
    .out   (_delay_fixed_32_0_1_108_2770_out)
  );
  delay_fixed_32_0_1_1727 delay_fixed_32_0_1_1727_2771 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2789:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4379),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1727_2771_out)
  );
  delay_fixed_32_0_1_207 delay_fixed_32_0_1_207_2772 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2790:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1816__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1962:116
    .out   (_delay_fixed_32_0_1_207_2772_out)
  );
  delay_fixed_32_0_1_249 delay_fixed_32_0_1_249_2773 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2791:146
    .clock (clock),
    .reset (reset),
    .in    (_dup689__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:835:111
    .out   (_delay_fixed_32_0_1_249_2773_out)
  );
  delay_fixed_1_0_0_79 delay_fixed_1_0_0_79_2774 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2792:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1823__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1969:139
    .out   (_delay_fixed_1_0_0_79_2774_out)
  );
  delay_fixed_32_0_1_1808 delay_fixed_32_0_1_1808_2775 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2793:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4361),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1808_2775_out)
  );
  delay_fixed_32_0_1_1659 delay_fixed_32_0_1_1659_2776 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2794:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4357),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1659_2776_out)
  );
  delay_fixed_32_0_1_65 delay_fixed_32_0_1_65_2777 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2795:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1820__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1966:154
    .out   (_delay_fixed_32_0_1_65_2777_out)
  );
  delay_fixed_32_0_1_1758 delay_fixed_32_0_1_1758_2778 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2796:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4361),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1758_2778_out)
  );
  delay_fixed_32_0_1_1693 delay_fixed_32_0_1_1693_2779 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2797:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4357),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1693_2779_out)
  );
  delay_fixed_32_0_1_65 delay_fixed_32_0_1_65_2780 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2798:142
    .clock (clock),
    .reset (reset),
    .in    (_dup684__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:830:111
    .out   (_delay_fixed_32_0_1_65_2780_out)
  );
  delay_fixed_32_0_1_207 delay_fixed_32_0_1_207_2781 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2799:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1816__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1962:116
    .out   (_delay_fixed_32_0_1_207_2781_out)
  );
  delay_fixed_32_0_1_90 delay_fixed_32_0_1_90_2782 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2800:142
    .clock (clock),
    .reset (reset),
    .in    (_dup680__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:826:111
    .out   (_delay_fixed_32_0_1_90_2782_out)
  );
  delay_fixed_1_0_0_18 delay_fixed_1_0_0_18_2783 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2801:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1813__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1959:139
    .out   (_delay_fixed_1_0_0_18_2783_out)
  );
  delay_fixed_32_0_1_1912 delay_fixed_32_0_1_1912_2784 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2802:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4339),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1912_2784_out)
  );
  delay_fixed_32_0_1_1826 delay_fixed_32_0_1_1826_2785 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2803:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4335),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1826_2785_out)
  );
  delay_fixed_32_0_1_58 delay_fixed_32_0_1_58_2786 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2804:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1810__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1956:154
    .out   (_delay_fixed_32_0_1_58_2786_out)
  );
  delay_fixed_32_0_1_1918 delay_fixed_32_0_1_1918_2787 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2805:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4339),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1918_2787_out)
  );
  delay_fixed_32_0_1_1860 delay_fixed_32_0_1_1860_2788 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2806:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4335),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1860_2788_out)
  );
  delay_fixed_32_0_1_537 delay_fixed_32_0_1_537_2789 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2807:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_1613),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_537_2789_out)
  );
  delay_fixed_32_0_1_442 delay_fixed_32_0_1_442_2790 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2808:146
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_1609),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_442_2790_out)
  );
  delay_fixed_32_0_1_98 delay_fixed_32_0_1_98_2791 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2809:142
    .clock (clock),
    .reset (reset),
    .in    (_dup670__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:816:111
    .out   (_delay_fixed_32_0_1_98_2791_out)
  );
  delay_fixed_32_0_1_445 delay_fixed_32_0_1_445_2792 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2810:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1806__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1952:116
    .out   (_delay_fixed_32_0_1_445_2792_out)
  );
  delay_fixed_32_0_1_584 delay_fixed_32_0_1_584_2793 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2811:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_1601),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_584_2793_out)
  );
  delay_fixed_32_0_1_417 delay_fixed_32_0_1_417_2794 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2812:146
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_1597),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_417_2794_out)
  );
  delay_fixed_32_0_1_98 delay_fixed_32_0_1_98_2795 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2813:142
    .clock (clock),
    .reset (reset),
    .in    (_dup670__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:816:111
    .out   (_delay_fixed_32_0_1_98_2795_out)
  );
  delay_fixed_32_0_1_19 delay_fixed_32_0_1_19_2796 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2814:142
    .clock (clock),
    .reset (reset),
    .in    (_MUX1802__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1948:169
    .out   (_delay_fixed_32_0_1_19_2796_out)
  );
  delay_fixed_32_0_1_1956 delay_fixed_32_0_1_1956_2797 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2815:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4317),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1956_2797_out)
  );
  delay_fixed_32_0_1_1874 delay_fixed_32_0_1_1874_2798 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2816:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4313),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1874_2798_out)
  );
  delay_fixed_32_0_1_51 delay_fixed_32_0_1_51_2799 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2817:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1800__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1946:154
    .out   (_delay_fixed_32_0_1_51_2799_out)
  );
  delay_fixed_32_0_1_1959 delay_fixed_32_0_1_1959_2800 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2818:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4317),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1959_2800_out)
  );
  delay_fixed_32_0_1_177 delay_fixed_32_0_1_177_2801 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2819:146
    .clock (clock),
    .reset (reset),
    .in    (_dup665__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:811:111
    .out   (_delay_fixed_32_0_1_177_2801_out)
  );
  delay_fixed_32_0_1_1908 delay_fixed_32_0_1_1908_2802 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2820:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4313),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1908_2802_out)
  );
  delay_fixed_32_0_1_177 delay_fixed_32_0_1_177_2803 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2821:146
    .clock (clock),
    .reset (reset),
    .in    (_dup665__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:811:111
    .out   (_delay_fixed_32_0_1_177_2803_out)
  );
  delay_fixed_32_0_1_440 delay_fixed_32_0_1_440_2804 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2822:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1796__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1942:116
    .out   (_delay_fixed_32_0_1_440_2804_out)
  );
  delay_fixed_32_0_1_258 delay_fixed_32_0_1_258_2805 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2823:146
    .clock (clock),
    .reset (reset),
    .in    (_dup661__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:807:111
    .out   (_delay_fixed_32_0_1_258_2805_out)
  );
  delay_fixed_32_0_1_258 delay_fixed_32_0_1_258_2806 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2824:146
    .clock (clock),
    .reset (reset),
    .in    (_dup661__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:807:111
    .out   (_delay_fixed_32_0_1_258_2806_out)
  );
  delay_fixed_1_0_0_53 delay_fixed_1_0_0_53_2807 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2825:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1793__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1939:139
    .out   (_delay_fixed_1_0_0_53_2807_out)
  );
  delay_fixed_32_0_1_1657 delay_fixed_32_0_1_1657_2808 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2826:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4295),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1657_2808_out)
  );
  delay_fixed_32_0_1_7 delay_fixed_32_0_1_7_2809 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2827:138
    .clock (clock),
    .reset (reset),
    .in    (_dup658__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:804:111
    .out   (_delay_fixed_32_0_1_7_2809_out)
  );
  delay_fixed_32_0_1_1542 delay_fixed_32_0_1_1542_2810 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2828:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4291),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1542_2810_out)
  );
  delay_fixed_32_0_1_7 delay_fixed_32_0_1_7_2811 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2829:138
    .clock (clock),
    .reset (reset),
    .in    (_dup658__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:804:111
    .out   (_delay_fixed_32_0_1_7_2811_out)
  );
  delay_fixed_32_0_1_57 delay_fixed_32_0_1_57_2812 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2830:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1790__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1936:154
    .out   (_delay_fixed_32_0_1_57_2812_out)
  );
  delay_fixed_32_0_1_1633 delay_fixed_32_0_1_1633_2813 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2831:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4295),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1633_2813_out)
  );
  delay_fixed_32_0_1_1576 delay_fixed_32_0_1_1576_2814 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2832:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4291),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1576_2814_out)
  );
  delay_fixed_32_0_1_30 delay_fixed_32_0_1_30_2815 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2833:142
    .clock (clock),
    .reset (reset),
    .in    (_dup653__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:799:111
    .out   (_delay_fixed_32_0_1_30_2815_out)
  );
  delay_fixed_32_0_1_30 delay_fixed_32_0_1_30_2816 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2834:142
    .clock (clock),
    .reset (reset),
    .in    (_dup653__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:799:111
    .out   (_delay_fixed_32_0_1_30_2816_out)
  );
  delay_fixed_32_0_1_158 delay_fixed_32_0_1_158_2817 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2835:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1786__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1932:116
    .out   (_delay_fixed_32_0_1_158_2817_out)
  );
  delay_fixed_32_0_1_132 delay_fixed_32_0_1_132_2818 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2836:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL651__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:797:131
    .out   (_delay_fixed_32_0_1_132_2818_out)
  );
  delay_fixed_32_0_1_186 delay_fixed_32_0_1_186_2819 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2837:146
    .clock (clock),
    .reset (reset),
    .in    (_dup49_const_fix_32_0_1__0000000000000235_1494),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
    .out   (_delay_fixed_32_0_1_186_2819_out)
  );
  delay_fixed_32_0_1_1685 delay_fixed_32_0_1_1685_2820 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2838:150
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_4280),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_1685_2820_out)
  );
  delay_fixed_32_0_1_247 delay_fixed_32_0_1_247_2821 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2839:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL648__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:794:131
    .out   (_delay_fixed_32_0_1_247_2821_out)
  );
  delay_fixed_32_0_1_1568 delay_fixed_32_0_1_1568_2822 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2840:150
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_4276),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_1568_2822_out)
  );
  delay_fixed_32_0_1_59 delay_fixed_32_0_1_59_2823 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2841:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1777__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1923:116
    .out   (_delay_fixed_32_0_1_59_2823_out)
  );
  delay_fixed_32_0_1_1 delay_fixed_32_0_1_1_2824 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2842:138
    .clock (clock),
    .reset (reset),
    .in    (_dup45_const_fix_32_0_1__0000000000000235_1494),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
    .out   (_delay_fixed_32_0_1_1_2824_out)
  );
  delay_fixed_32_0_1_229 delay_fixed_32_0_1_229_2825 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2843:146
    .clock (clock),
    .reset (reset),
    .in    (_dup43_const_fix_32_0_1__0000000000000235_1494),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
    .out   (_delay_fixed_32_0_1_229_2825_out)
  );
  delay_fixed_32_0_1_1646 delay_fixed_32_0_1_1646_2826 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2844:150
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_4268),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_1646_2826_out)
  );
  delay_fixed_32_0_1_129 delay_fixed_32_0_1_129_2827 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2845:146
    .clock (clock),
    .reset (reset),
    .in    (_dup645__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:791:111
    .out   (_delay_fixed_32_0_1_129_2827_out)
  );
  delay_fixed_32_0_1_1500 delay_fixed_32_0_1_1500_2828 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2846:150
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_4264),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_1500_2828_out)
  );
  delay_fixed_32_0_1_59 delay_fixed_32_0_1_59_2829 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2847:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1777__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1923:116
    .out   (_delay_fixed_32_0_1_59_2829_out)
  );
  delay_fixed_32_0_1_2 delay_fixed_32_0_1_2_2830 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2848:138
    .clock (clock),
    .reset (reset),
    .in    (_dup641__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:787:111
    .out   (_delay_fixed_32_0_1_2_2830_out)
  );
  delay_fixed_32_0_1_2 delay_fixed_32_0_1_2_2831 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2849:138
    .clock (clock),
    .reset (reset),
    .in    (_dup641__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:787:111
    .out   (_delay_fixed_32_0_1_2_2831_out)
  );
  delay_fixed_32_0_1_76 delay_fixed_32_0_1_76_2832 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2850:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1772__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1918:116
    .out   (_delay_fixed_32_0_1_76_2832_out)
  );
  delay_fixed_32_0_1_76 delay_fixed_32_0_1_76_2833 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2851:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1772__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1918:116
    .out   (_delay_fixed_32_0_1_76_2833_out)
  );
  delay_fixed_32_0_1_11 delay_fixed_32_0_1_11_2834 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2852:142
    .clock (clock),
    .reset (reset),
    .in    (_dup636__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:782:111
    .out   (_delay_fixed_32_0_1_11_2834_out)
  );
  delay_fixed_32_0_1_127 delay_fixed_32_0_1_127_2835 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2853:146
    .clock (clock),
    .reset (reset),
    .in    (_dup33_const_fix_32_0_1__0000000000000235_1494),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
    .out   (_delay_fixed_32_0_1_127_2835_out)
  );
  delay_fixed_32_0_1_70 delay_fixed_32_0_1_70_2836 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2854:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1768__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1914:116
    .out   (_delay_fixed_32_0_1_70_2836_out)
  );
  delay_fixed_32_0_1_61 delay_fixed_32_0_1_61_2837 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2855:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL635__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:781:131
    .out   (_delay_fixed_32_0_1_61_2837_out)
  );
  delay_fixed_32_0_1_70 delay_fixed_32_0_1_70_2838 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2856:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1768__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1914:116
    .out   (_delay_fixed_32_0_1_70_2838_out)
  );
  delay_fixed_32_0_1_40 delay_fixed_32_0_1_40_2839 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2857:142
    .clock (clock),
    .reset (reset),
    .in    (_dup29_const_fix_32_0_1__0000000000000235_1494),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
    .out   (_delay_fixed_32_0_1_40_2839_out)
  );
  delay_fixed_32_0_1_164 delay_fixed_32_0_1_164_2840 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2858:146
    .clock (clock),
    .reset (reset),
    .in    (_dup27_const_fix_32_0_1__0000000000000235_1494),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
    .out   (_delay_fixed_32_0_1_164_2840_out)
  );
  delay_fixed_32_0_1_7 delay_fixed_32_0_1_7_2841 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2859:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1764__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1910:116
    .out   (_delay_fixed_32_0_1_7_2841_out)
  );
  delay_fixed_32_0_1_29 delay_fixed_32_0_1_29_2842 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2860:142
    .clock (clock),
    .reset (reset),
    .in    (_dup631__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:777:111
    .out   (_delay_fixed_32_0_1_29_2842_out)
  );
  delay_fixed_32_0_1_7 delay_fixed_32_0_1_7_2843 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2861:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1764__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1910:116
    .out   (_delay_fixed_32_0_1_7_2843_out)
  );
  delay_fixed_32_0_1_30 delay_fixed_32_0_1_30_2844 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2862:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL629__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:775:131
    .out   (_delay_fixed_32_0_1_30_2844_out)
  );
  delay_fixed_32_0_1_38 delay_fixed_32_0_1_38_2845 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2863:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1761__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1907:116
    .out   (_delay_fixed_32_0_1_38_2845_out)
  );
  delay_fixed_32_0_1_146 delay_fixed_32_0_1_146_2846 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2864:146
    .clock (clock),
    .reset (reset),
    .in    (_dup21_const_fix_32_0_1__0000000000000235_1494),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
    .out   (_delay_fixed_32_0_1_146_2846_out)
  );
  delay_fixed_32_0_1_38 delay_fixed_32_0_1_38_2847 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2865:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1761__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1907:116
    .out   (_delay_fixed_32_0_1_38_2847_out)
  );
  delay_fixed_32_0_1_24 delay_fixed_32_0_1_24_2848 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2866:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL626__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:772:131
    .out   (_delay_fixed_32_0_1_24_2848_out)
  );
  delay_fixed_32_0_1_175 delay_fixed_32_0_1_175_2849 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2867:146
    .clock (clock),
    .reset (reset),
    .in    (_dup17_const_fix_32_0_1__0000000000000235_1494),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
    .out   (_delay_fixed_32_0_1_175_2849_out)
  );
  delay_fixed_32_0_1_202 delay_fixed_32_0_1_202_2850 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2868:146
    .clock (clock),
    .reset (reset),
    .in    (_dup15_const_fix_32_0_1__0000000000000235_1494),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
    .out   (_delay_fixed_32_0_1_202_2850_out)
  );
  delay_fixed_32_0_1_130 delay_fixed_32_0_1_130_2851 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2869:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1757__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1903:136
    .out   (_delay_fixed_32_0_1_130_2851_out)
  );
  delay_fixed_32_0_1_73 delay_fixed_32_0_1_73_2852 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2870:142
    .clock (clock),
    .reset (reset),
    .in    (_dup623__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:769:111
    .out   (_delay_fixed_32_0_1_73_2852_out)
  );
  delay_fixed_32_0_1_113 delay_fixed_32_0_1_113_2853 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2871:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_1488),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_113_2853_out)
  );
  delay_fixed_32_0_1_35 delay_fixed_32_0_1_35_2854 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2872:142
    .clock (clock),
    .reset (reset),
    .in    (_dup579__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:725:111
    .out   (_delay_fixed_32_0_1_35_2854_out)
  );
  delay_fixed_32_0_1_134 delay_fixed_32_0_1_134_2855 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2873:146
    .clock (clock),
    .reset (reset),
    .in    (_dup584__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:730:111
    .out   (_delay_fixed_32_0_1_134_2855_out)
  );
  delay_fixed_32_0_1_198 delay_fixed_32_0_1_198_2856 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2874:146
    .clock (clock),
    .reset (reset),
    .in    (_dup589__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:735:111
    .out   (_delay_fixed_32_0_1_198_2856_out)
  );
  delay_fixed_32_0_1_73 delay_fixed_32_0_1_73_2857 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2875:142
    .clock (clock),
    .reset (reset),
    .in    (_dup595__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:741:111
    .out   (_delay_fixed_32_0_1_73_2857_out)
  );
  delay_fixed_32_0_1_73 delay_fixed_32_0_1_73_2858 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2876:142
    .clock (clock),
    .reset (reset),
    .in    (_dup595__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:741:111
    .out   (_delay_fixed_32_0_1_73_2858_out)
  );
  delay_fixed_32_0_1_198 delay_fixed_32_0_1_198_2859 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2877:146
    .clock (clock),
    .reset (reset),
    .in    (_dup589__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:735:111
    .out   (_delay_fixed_32_0_1_198_2859_out)
  );
  delay_fixed_32_0_1_134 delay_fixed_32_0_1_134_2860 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2878:146
    .clock (clock),
    .reset (reset),
    .in    (_dup584__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:730:111
    .out   (_delay_fixed_32_0_1_134_2860_out)
  );
  delay_fixed_32_0_1_35 delay_fixed_32_0_1_35_2861 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2879:142
    .clock (clock),
    .reset (reset),
    .in    (_dup579__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:725:111
    .out   (_delay_fixed_32_0_1_35_2861_out)
  );
  delay_fixed_32_0_1_670 delay_fixed_32_0_1_670_2862 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2880:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_1382),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_670_2862_out)
  );
  delay_fixed_32_0_1_516 delay_fixed_32_0_1_516_2863 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2881:146
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_1378),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_516_2863_out)
  );
  delay_fixed_32_0_1_94 delay_fixed_32_0_1_94_2864 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2882:142
    .clock (clock),
    .reset (reset),
    .in    (_dup569__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:715:111
    .out   (_delay_fixed_32_0_1_94_2864_out)
  );
  delay_fixed_32_0_1_610 delay_fixed_32_0_1_610_2865 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2883:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_1370),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_610_2865_out)
  );
  delay_fixed_32_0_1_497 delay_fixed_32_0_1_497_2866 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2884:146
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_1366),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_497_2866_out)
  );
  delay_fixed_32_0_1_94 delay_fixed_32_0_1_94_2867 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2885:142
    .clock (clock),
    .reset (reset),
    .in    (_dup569__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:715:111
    .out   (_delay_fixed_32_0_1_94_2867_out)
  );
  delay_fixed_32_0_1_174 delay_fixed_32_0_1_174_2868 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2886:146
    .clock (clock),
    .reset (reset),
    .in    (_dup565__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:711:111
    .out   (_delay_fixed_32_0_1_174_2868_out)
  );
  delay_fixed_32_0_1_174 delay_fixed_32_0_1_174_2869 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2887:146
    .clock (clock),
    .reset (reset),
    .in    (_dup565__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:711:111
    .out   (_delay_fixed_32_0_1_174_2869_out)
  );
  delay_fixed_32_0_1_118 delay_fixed_32_0_1_118_2870 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2888:146
    .clock (clock),
    .reset (reset),
    .in    (_dup561__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:707:111
    .out   (_delay_fixed_32_0_1_118_2870_out)
  );
  delay_fixed_32_0_1_118 delay_fixed_32_0_1_118_2871 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2889:146
    .clock (clock),
    .reset (reset),
    .in    (_dup561__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:707:111
    .out   (_delay_fixed_32_0_1_118_2871_out)
  );
  delay_fixed_32_0_1_57 delay_fixed_32_0_1_57_2872 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2890:142
    .clock (clock),
    .reset (reset),
    .in    (_dup558__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:704:111
    .out   (_delay_fixed_32_0_1_57_2872_out)
  );
  delay_fixed_32_0_1_57 delay_fixed_32_0_1_57_2873 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2891:142
    .clock (clock),
    .reset (reset),
    .in    (_dup558__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:704:111
    .out   (_delay_fixed_32_0_1_57_2873_out)
  );
  delay_fixed_32_0_1_1 delay_fixed_32_0_1_1_2874 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2892:138
    .clock (clock),
    .reset (reset),
    .in    (_dup553__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:699:111
    .out   (_delay_fixed_32_0_1_1_2874_out)
  );
  delay_fixed_32_0_1_1 delay_fixed_32_0_1_1_2875 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2893:138
    .clock (clock),
    .reset (reset),
    .in    (_dup553__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:699:111
    .out   (_delay_fixed_32_0_1_1_2875_out)
  );
  delay_fixed_32_0_1_95 delay_fixed_32_0_1_95_2876 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2894:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL551__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:697:131
    .out   (_delay_fixed_32_0_1_95_2876_out)
  );
  delay_fixed_32_0_1_122 delay_fixed_32_0_1_122_2877 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2895:146
    .clock (clock),
    .reset (reset),
    .in    (_dup49_const_fix_32_0_1__0000000000000235_1263),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
    .out   (_delay_fixed_32_0_1_122_2877_out)
  );
  delay_fixed_32_0_1_110 delay_fixed_32_0_1_110_2878 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2896:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL548__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:694:131
    .out   (_delay_fixed_32_0_1_110_2878_out)
  );
  delay_fixed_32_0_1_64 delay_fixed_32_0_1_64_2879 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2897:142
    .clock (clock),
    .reset (reset),
    .in    (_dup45_const_fix_32_0_1__0000000000000235_1263),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
    .out   (_delay_fixed_32_0_1_64_2879_out)
  );
  delay_fixed_32_0_1_177 delay_fixed_32_0_1_177_2880 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2898:146
    .clock (clock),
    .reset (reset),
    .in    (_dup43_const_fix_32_0_1__0000000000000235_1263),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
    .out   (_delay_fixed_32_0_1_177_2880_out)
  );
  delay_fixed_32_0_1_2 delay_fixed_32_0_1_2_2881 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2899:138
    .clock (clock),
    .reset (reset),
    .in    (_dup545__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:691:111
    .out   (_delay_fixed_32_0_1_2_2881_out)
  );
  delay_fixed_32_0_1_23 delay_fixed_32_0_1_23_2882 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2900:142
    .clock (clock),
    .reset (reset),
    .in    (_dup541__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:687:111
    .out   (_delay_fixed_32_0_1_23_2882_out)
  );
  delay_fixed_32_0_1_23 delay_fixed_32_0_1_23_2883 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2901:142
    .clock (clock),
    .reset (reset),
    .in    (_dup541__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:687:111
    .out   (_delay_fixed_32_0_1_23_2883_out)
  );
  delay_fixed_32_0_1_3 delay_fixed_32_0_1_3_2884 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2902:138
    .clock (clock),
    .reset (reset),
    .in    (_dup536__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:682:111
    .out   (_delay_fixed_32_0_1_3_2884_out)
  );
  delay_fixed_32_0_1_138 delay_fixed_32_0_1_138_2885 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2903:146
    .clock (clock),
    .reset (reset),
    .in    (_dup33_const_fix_32_0_1__0000000000000235_1263),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
    .out   (_delay_fixed_32_0_1_138_2885_out)
  );
  delay_fixed_32_0_1_103 delay_fixed_32_0_1_103_2886 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2904:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL535__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:681:131
    .out   (_delay_fixed_32_0_1_103_2886_out)
  );
  delay_fixed_32_0_1_10 delay_fixed_32_0_1_10_2887 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2905:142
    .clock (clock),
    .reset (reset),
    .in    (_dup29_const_fix_32_0_1__0000000000000235_1263),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
    .out   (_delay_fixed_32_0_1_10_2887_out)
  );
  delay_fixed_32_0_1_145 delay_fixed_32_0_1_145_2888 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2906:146
    .clock (clock),
    .reset (reset),
    .in    (_dup27_const_fix_32_0_1__0000000000000235_1263),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
    .out   (_delay_fixed_32_0_1_145_2888_out)
  );
  delay_fixed_32_0_1_70 delay_fixed_32_0_1_70_2889 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2907:142
    .clock (clock),
    .reset (reset),
    .in    (_dup531__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:677:111
    .out   (_delay_fixed_32_0_1_70_2889_out)
  );
  delay_fixed_32_0_1_131 delay_fixed_32_0_1_131_2890 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2908:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL529__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:675:131
    .out   (_delay_fixed_32_0_1_131_2890_out)
  );
  delay_fixed_32_0_1_57 delay_fixed_32_0_1_57_2891 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2909:142
    .clock (clock),
    .reset (reset),
    .in    (_dup479__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:625:111
    .out   (_delay_fixed_32_0_1_57_2891_out)
  );
  delay_fixed_32_0_1_272 delay_fixed_32_0_1_272_2892 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2910:146
    .clock (clock),
    .reset (reset),
    .in    (_dup484__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:630:111
    .out   (_delay_fixed_32_0_1_272_2892_out)
  );
  delay_fixed_32_0_1_212 delay_fixed_32_0_1_212_2893 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2911:146
    .clock (clock),
    .reset (reset),
    .in    (_dup489__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:635:111
    .out   (_delay_fixed_32_0_1_212_2893_out)
  );
  delay_fixed_32_0_1_37 delay_fixed_32_0_1_37_2894 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2912:142
    .clock (clock),
    .reset (reset),
    .in    (_dup495__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:641:111
    .out   (_delay_fixed_32_0_1_37_2894_out)
  );
  delay_fixed_32_0_1_37 delay_fixed_32_0_1_37_2895 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2913:142
    .clock (clock),
    .reset (reset),
    .in    (_dup495__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:641:111
    .out   (_delay_fixed_32_0_1_37_2895_out)
  );
  delay_fixed_32_0_1_212 delay_fixed_32_0_1_212_2896 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2914:146
    .clock (clock),
    .reset (reset),
    .in    (_dup489__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:635:111
    .out   (_delay_fixed_32_0_1_212_2896_out)
  );
  delay_fixed_32_0_1_272 delay_fixed_32_0_1_272_2897 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2915:146
    .clock (clock),
    .reset (reset),
    .in    (_dup484__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:630:111
    .out   (_delay_fixed_32_0_1_272_2897_out)
  );
  delay_fixed_32_0_1_57 delay_fixed_32_0_1_57_2898 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2916:142
    .clock (clock),
    .reset (reset),
    .in    (_dup479__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:625:111
    .out   (_delay_fixed_32_0_1_57_2898_out)
  );
  delay_fixed_32_0_1_561 delay_fixed_32_0_1_561_2899 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2917:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_1151),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_561_2899_out)
  );
  delay_fixed_32_0_1_473 delay_fixed_32_0_1_473_2900 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2918:146
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_1147),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_473_2900_out)
  );
  delay_fixed_32_0_1_103 delay_fixed_32_0_1_103_2901 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2919:146
    .clock (clock),
    .reset (reset),
    .in    (_dup470__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:616:111
    .out   (_delay_fixed_32_0_1_103_2901_out)
  );
  delay_fixed_32_0_1_605 delay_fixed_32_0_1_605_2902 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2920:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_1139),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_605_2902_out)
  );
  delay_fixed_32_0_1_504 delay_fixed_32_0_1_504_2903 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2921:146
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_1135),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_504_2903_out)
  );
  delay_fixed_32_0_1_103 delay_fixed_32_0_1_103_2904 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2922:146
    .clock (clock),
    .reset (reset),
    .in    (_dup470__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:616:111
    .out   (_delay_fixed_32_0_1_103_2904_out)
  );
  delay_fixed_32_0_1_47 delay_fixed_32_0_1_47_2905 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2923:142
    .clock (clock),
    .reset (reset),
    .in    (_dup466__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:612:111
    .out   (_delay_fixed_32_0_1_47_2905_out)
  );
  delay_fixed_32_0_1_47 delay_fixed_32_0_1_47_2906 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2924:142
    .clock (clock),
    .reset (reset),
    .in    (_dup466__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:612:111
    .out   (_delay_fixed_32_0_1_47_2906_out)
  );
  delay_fixed_32_0_1_45 delay_fixed_32_0_1_45_2907 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2925:142
    .clock (clock),
    .reset (reset),
    .in    (_dup461__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:607:111
    .out   (_delay_fixed_32_0_1_45_2907_out)
  );
  delay_fixed_32_0_1_45 delay_fixed_32_0_1_45_2908 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2926:142
    .clock (clock),
    .reset (reset),
    .in    (_dup461__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:607:111
    .out   (_delay_fixed_32_0_1_45_2908_out)
  );
  delay_fixed_32_0_1_40 delay_fixed_32_0_1_40_2909 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2927:142
    .clock (clock),
    .reset (reset),
    .in    (_dup457__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:603:111
    .out   (_delay_fixed_32_0_1_40_2909_out)
  );
  delay_fixed_32_0_1_40 delay_fixed_32_0_1_40_2910 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2928:142
    .clock (clock),
    .reset (reset),
    .in    (_dup457__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:603:111
    .out   (_delay_fixed_32_0_1_40_2910_out)
  );
  delay_fixed_32_0_1_72 delay_fixed_32_0_1_72_2911 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2929:142
    .clock (clock),
    .reset (reset),
    .in    (_dup453__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:599:111
    .out   (_delay_fixed_32_0_1_72_2911_out)
  );
  delay_fixed_32_0_1_72 delay_fixed_32_0_1_72_2912 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2930:142
    .clock (clock),
    .reset (reset),
    .in    (_dup453__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:599:111
    .out   (_delay_fixed_32_0_1_72_2912_out)
  );
  delay_fixed_32_0_1_163 delay_fixed_32_0_1_163_2913 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2931:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL451__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:597:131
    .out   (_delay_fixed_32_0_1_163_2913_out)
  );
  delay_fixed_32_0_1_71 delay_fixed_32_0_1_71_2914 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2932:142
    .clock (clock),
    .reset (reset),
    .in    (_dup49_const_fix_32_0_1__0000000000000235_1032),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
    .out   (_delay_fixed_32_0_1_71_2914_out)
  );
  delay_fixed_32_0_1_76 delay_fixed_32_0_1_76_2915 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2933:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL448__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:594:131
    .out   (_delay_fixed_32_0_1_76_2915_out)
  );
  delay_fixed_32_0_1_81 delay_fixed_32_0_1_81_2916 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2934:142
    .clock (clock),
    .reset (reset),
    .in    (_dup45_const_fix_32_0_1__0000000000000235_1032),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
    .out   (_delay_fixed_32_0_1_81_2916_out)
  );
  delay_fixed_32_0_1_131 delay_fixed_32_0_1_131_2917 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2935:146
    .clock (clock),
    .reset (reset),
    .in    (_dup43_const_fix_32_0_1__0000000000000235_1032),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
    .out   (_delay_fixed_32_0_1_131_2917_out)
  );
  delay_fixed_32_0_1_66 delay_fixed_32_0_1_66_2918 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2936:142
    .clock (clock),
    .reset (reset),
    .in    (_dup444__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:590:111
    .out   (_delay_fixed_32_0_1_66_2918_out)
  );
  delay_fixed_32_0_1_4 delay_fixed_32_0_1_4_2919 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2937:138
    .clock (clock),
    .reset (reset),
    .in    (_dup441__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:587:111
    .out   (_delay_fixed_32_0_1_4_2919_out)
  );
  delay_fixed_32_0_1_4 delay_fixed_32_0_1_4_2920 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2938:138
    .clock (clock),
    .reset (reset),
    .in    (_dup441__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:587:111
    .out   (_delay_fixed_32_0_1_4_2920_out)
  );
  delay_fixed_32_0_1_166 delay_fixed_32_0_1_166_2921 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2939:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL438__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:584:131
    .out   (_delay_fixed_32_0_1_166_2921_out)
  );
  delay_fixed_32_0_1_79 delay_fixed_32_0_1_79_2922 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2940:142
    .clock (clock),
    .reset (reset),
    .in    (_dup33_const_fix_32_0_1__0000000000000235_1032),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
    .out   (_delay_fixed_32_0_1_79_2922_out)
  );
  delay_fixed_32_0_1_150 delay_fixed_32_0_1_150_2923 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2941:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL435__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:581:131
    .out   (_delay_fixed_32_0_1_150_2923_out)
  );
  delay_fixed_32_0_1_10 delay_fixed_32_0_1_10_2924 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2942:142
    .clock (clock),
    .reset (reset),
    .in    (_dup29_const_fix_32_0_1__0000000000000235_1032),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
    .out   (_delay_fixed_32_0_1_10_2924_out)
  );
  delay_fixed_32_0_1_114 delay_fixed_32_0_1_114_2925 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2943:146
    .clock (clock),
    .reset (reset),
    .in    (_dup27_const_fix_32_0_1__0000000000000235_1032),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
    .out   (_delay_fixed_32_0_1_114_2925_out)
  );
  delay_fixed_32_0_1_11 delay_fixed_32_0_1_11_2926 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2944:142
    .clock (clock),
    .reset (reset),
    .in    (_dup431__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:577:111
    .out   (_delay_fixed_32_0_1_11_2926_out)
  );
  delay_fixed_32_0_1_89 delay_fixed_32_0_1_89_2927 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2945:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL429__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:575:131
    .out   (_delay_fixed_32_0_1_89_2927_out)
  );
  delay_fixed_32_0_1_21 delay_fixed_32_0_1_21_2928 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2946:142
    .clock (clock),
    .reset (reset),
    .in    (_dup21_const_fix_32_0_1__0000000000000235_1032),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
    .out   (_delay_fixed_32_0_1_21_2928_out)
  );
  delay_fixed_32_0_1_31 delay_fixed_32_0_1_31_2929 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2947:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL426__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:572:131
    .out   (_delay_fixed_32_0_1_31_2929_out)
  );
  delay_fixed_32_0_1_7 delay_fixed_32_0_1_7_2930 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2948:138
    .clock (clock),
    .reset (reset),
    .in    (_dup17_const_fix_32_0_1__0000000000000235_1032),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
    .out   (_delay_fixed_32_0_1_7_2930_out)
  );
  delay_fixed_32_0_1_91 delay_fixed_32_0_1_91_2931 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2949:142
    .clock (clock),
    .reset (reset),
    .in    (_dup15_const_fix_32_0_1__0000000000000235_1032),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
    .out   (_delay_fixed_32_0_1_91_2931_out)
  );
  delay_fixed_32_0_1_30 delay_fixed_32_0_1_30_2932 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2950:142
    .clock (clock),
    .reset (reset),
    .in    (_dup423__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:569:111
    .out   (_delay_fixed_32_0_1_30_2932_out)
  );
  delay_fixed_32_0_1_109 delay_fixed_32_0_1_109_2933 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2951:146
    .clock (clock),
    .reset (reset),
    .in    (_dup21_const_fix_32_0_1__0000000000000235_1263),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
    .out   (_delay_fixed_32_0_1_109_2933_out)
  );
  delay_fixed_32_0_1_166 delay_fixed_32_0_1_166_2934 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2952:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_1026),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_166_2934_out)
  );
  delay_fixed_32_0_1_57 delay_fixed_32_0_1_57_2935 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2953:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL526__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:672:131
    .out   (_delay_fixed_32_0_1_57_2935_out)
  );
  delay_fixed_32_0_1_75 delay_fixed_32_0_1_75_2936 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2954:142
    .clock (clock),
    .reset (reset),
    .in    (_dup17_const_fix_32_0_1__0000000000000235_1263),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
    .out   (_delay_fixed_32_0_1_75_2936_out)
  );
  delay_fixed_32_0_1_162 delay_fixed_32_0_1_162_2937 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2955:146
    .clock (clock),
    .reset (reset),
    .in    (_dup15_const_fix_32_0_1__0000000000000235_1263),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
    .out   (_delay_fixed_32_0_1_162_2937_out)
  );
  delay_fixed_32_0_1_10 delay_fixed_32_0_1_10_2938 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2956:142
    .clock (clock),
    .reset (reset),
    .in    (_dup523__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:669:111
    .out   (_delay_fixed_32_0_1_10_2938_out)
  );
  delay_fixed_32_0_1_132 delay_fixed_32_0_1_132_2939 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2957:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_1257),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_132_2939_out)
  );
  delay_fixed_32_0_1_55 delay_fixed_32_0_1_55_2940 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2958:142
    .clock (clock),
    .reset (reset),
    .in    (_dup380__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:526:111
    .out   (_delay_fixed_32_0_1_55_2940_out)
  );
  delay_fixed_32_0_1_270 delay_fixed_32_0_1_270_2941 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2959:146
    .clock (clock),
    .reset (reset),
    .in    (_dup384__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:530:111
    .out   (_delay_fixed_32_0_1_270_2941_out)
  );
  delay_fixed_32_0_1_55 delay_fixed_32_0_1_55_2942 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2960:142
    .clock (clock),
    .reset (reset),
    .in    (_dup380__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:526:111
    .out   (_delay_fixed_32_0_1_55_2942_out)
  );
  delay_fixed_32_0_1_609 delay_fixed_32_0_1_609_2943 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2961:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_920),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_609_2943_out)
  );
  delay_fixed_32_0_1_456 delay_fixed_32_0_1_456_2944 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2962:146
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_916),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_456_2944_out)
  );
  delay_fixed_32_0_1_46 delay_fixed_32_0_1_46_2945 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2963:142
    .clock (clock),
    .reset (reset),
    .in    (_dup370__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:516:111
    .out   (_delay_fixed_32_0_1_46_2945_out)
  );
  delay_fixed_32_0_1_625 delay_fixed_32_0_1_625_2946 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2964:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_908),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_625_2946_out)
  );
  delay_fixed_32_0_1_482 delay_fixed_32_0_1_482_2947 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2965:146
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_904),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_482_2947_out)
  );
  delay_fixed_32_0_1_46 delay_fixed_32_0_1_46_2948 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2966:142
    .clock (clock),
    .reset (reset),
    .in    (_dup370__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:516:111
    .out   (_delay_fixed_32_0_1_46_2948_out)
  );
  delay_fixed_32_0_1_87 delay_fixed_32_0_1_87_2949 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2967:142
    .clock (clock),
    .reset (reset),
    .in    (_dup365__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:511:111
    .out   (_delay_fixed_32_0_1_87_2949_out)
  );
  delay_fixed_32_0_1_87 delay_fixed_32_0_1_87_2950 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2968:142
    .clock (clock),
    .reset (reset),
    .in    (_dup365__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:511:111
    .out   (_delay_fixed_32_0_1_87_2950_out)
  );
  delay_fixed_32_0_1_14 delay_fixed_32_0_1_14_2951 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2969:142
    .clock (clock),
    .reset (reset),
    .in    (_dup361__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:507:111
    .out   (_delay_fixed_32_0_1_14_2951_out)
  );
  delay_fixed_32_0_1_14 delay_fixed_32_0_1_14_2952 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2970:142
    .clock (clock),
    .reset (reset),
    .in    (_dup361__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:507:111
    .out   (_delay_fixed_32_0_1_14_2952_out)
  );
  delay_fixed_32_0_1_16 delay_fixed_32_0_1_16_2953 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2971:142
    .clock (clock),
    .reset (reset),
    .in    (_dup357__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:503:111
    .out   (_delay_fixed_32_0_1_16_2953_out)
  );
  delay_fixed_32_0_1_16 delay_fixed_32_0_1_16_2954 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2972:142
    .clock (clock),
    .reset (reset),
    .in    (_dup357__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:503:111
    .out   (_delay_fixed_32_0_1_16_2954_out)
  );
  delay_fixed_32_0_1_15 delay_fixed_32_0_1_15_2955 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2973:142
    .clock (clock),
    .reset (reset),
    .in    (_dup353__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:499:111
    .out   (_delay_fixed_32_0_1_15_2955_out)
  );
  delay_fixed_32_0_1_15 delay_fixed_32_0_1_15_2956 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2974:142
    .clock (clock),
    .reset (reset),
    .in    (_dup353__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:499:111
    .out   (_delay_fixed_32_0_1_15_2956_out)
  );
  delay_fixed_32_0_1_253 delay_fixed_32_0_1_253_2957 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2975:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL351__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:497:131
    .out   (_delay_fixed_32_0_1_253_2957_out)
  );
  delay_fixed_32_0_1_28 delay_fixed_32_0_1_28_2958 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2976:142
    .clock (clock),
    .reset (reset),
    .in    (_dup49_const_fix_32_0_1__0000000000000235_801),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
    .out   (_delay_fixed_32_0_1_28_2958_out)
  );
  delay_fixed_32_0_1_155 delay_fixed_32_0_1_155_2959 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2977:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL348__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:494:131
    .out   (_delay_fixed_32_0_1_155_2959_out)
  );
  delay_fixed_32_0_1_44 delay_fixed_32_0_1_44_2960 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2978:142
    .clock (clock),
    .reset (reset),
    .in    (_dup45_const_fix_32_0_1__0000000000000235_801),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
    .out   (_delay_fixed_32_0_1_44_2960_out)
  );
  delay_fixed_32_0_1_136 delay_fixed_32_0_1_136_2961 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2979:146
    .clock (clock),
    .reset (reset),
    .in    (_dup43_const_fix_32_0_1__0000000000000235_801),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
    .out   (_delay_fixed_32_0_1_136_2961_out)
  );
  delay_fixed_32_0_1_72 delay_fixed_32_0_1_72_2962 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2980:142
    .clock (clock),
    .reset (reset),
    .in    (_dup344__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:490:111
    .out   (_delay_fixed_32_0_1_72_2962_out)
  );
  delay_fixed_32_0_1_12 delay_fixed_32_0_1_12_2963 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2981:142
    .clock (clock),
    .reset (reset),
    .in    (_dup340__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:486:111
    .out   (_delay_fixed_32_0_1_12_2963_out)
  );
  delay_fixed_32_0_1_12 delay_fixed_32_0_1_12_2964 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2982:142
    .clock (clock),
    .reset (reset),
    .in    (_dup340__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:486:111
    .out   (_delay_fixed_32_0_1_12_2964_out)
  );
  delay_fixed_32_0_1_186 delay_fixed_32_0_1_186_2965 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2983:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL338__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:484:131
    .out   (_delay_fixed_32_0_1_186_2965_out)
  );
  delay_fixed_32_0_1_25 delay_fixed_32_0_1_25_2966 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2984:142
    .clock (clock),
    .reset (reset),
    .in    (_dup33_const_fix_32_0_1__0000000000000235_801),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
    .out   (_delay_fixed_32_0_1_25_2966_out)
  );
  delay_fixed_32_0_1_94 delay_fixed_32_0_1_94_2967 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2985:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL335__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:481:131
    .out   (_delay_fixed_32_0_1_94_2967_out)
  );
  delay_fixed_32_0_1_43 delay_fixed_32_0_1_43_2968 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2986:142
    .clock (clock),
    .reset (reset),
    .in    (_dup29_const_fix_32_0_1__0000000000000235_801),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
    .out   (_delay_fixed_32_0_1_43_2968_out)
  );
  delay_fixed_32_0_1_199 delay_fixed_32_0_1_199_2969 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2987:146
    .clock (clock),
    .reset (reset),
    .in    (_dup27_const_fix_32_0_1__0000000000000235_801),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
    .out   (_delay_fixed_32_0_1_199_2969_out)
  );
  delay_fixed_32_0_1_76 delay_fixed_32_0_1_76_2970 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2988:142
    .clock (clock),
    .reset (reset),
    .in    (_dup332__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:478:111
    .out   (_delay_fixed_32_0_1_76_2970_out)
  );
  delay_fixed_32_0_1_39 delay_fixed_32_0_1_39_2971 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2989:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL329__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:475:131
    .out   (_delay_fixed_32_0_1_39_2971_out)
  );
  delay_fixed_32_0_1_142 delay_fixed_32_0_1_142_2972 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2990:146
    .clock (clock),
    .reset (reset),
    .in    (_dup21_const_fix_32_0_1__0000000000000235_801),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
    .out   (_delay_fixed_32_0_1_142_2972_out)
  );
  delay_fixed_32_0_1_60 delay_fixed_32_0_1_60_2973 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2991:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL326__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:472:131
    .out   (_delay_fixed_32_0_1_60_2973_out)
  );
  delay_fixed_32_0_1_44 delay_fixed_32_0_1_44_2974 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2992:142
    .clock (clock),
    .reset (reset),
    .in    (_dup17_const_fix_32_0_1__0000000000000235_801),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
    .out   (_delay_fixed_32_0_1_44_2974_out)
  );
  delay_fixed_32_0_1_113 delay_fixed_32_0_1_113_2975 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2993:146
    .clock (clock),
    .reset (reset),
    .in    (_dup15_const_fix_32_0_1__0000000000000235_801),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
    .out   (_delay_fixed_32_0_1_113_2975_out)
  );
  delay_fixed_32_0_1_54 delay_fixed_32_0_1_54_2976 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2994:142
    .clock (clock),
    .reset (reset),
    .in    (_dup322__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:468:111
    .out   (_delay_fixed_32_0_1_54_2976_out)
  );
  delay_fixed_32_0_1_122 delay_fixed_32_0_1_122_2977 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2995:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_795),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_122_2977_out)
  );
  delay_fixed_32_0_1_190 delay_fixed_32_0_1_190_2978 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2996:146
    .clock (clock),
    .reset (reset),
    .in    (_dup890__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1036:111
    .out   (_delay_fixed_32_0_1_190_2978_out)
  );
  delay_fixed_32_0_1_1564 delay_fixed_32_0_1_1564_2979 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2997:150
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_2096),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_1564_2979_out)
  );
  delay_fixed_32_0_1_1391 delay_fixed_32_0_1_1391_2980 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2998:150
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_2092),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_1391_2980_out)
  );
  delay_fixed_32_0_1_6 delay_fixed_32_0_1_6_2981 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2999:138
    .clock (clock),
    .reset (reset),
    .in    (_dup881__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1027:111
    .out   (_delay_fixed_32_0_1_6_2981_out)
  );
  delay_fixed_32_0_1_70 delay_fixed_32_0_1_70_2982 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3000:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1019__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1165:116
    .out   (_delay_fixed_32_0_1_70_2982_out)
  );
  delay_fixed_32_0_1_1557 delay_fixed_32_0_1_1557_2983 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3001:150
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_2084),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_1557_2983_out)
  );
  delay_fixed_32_0_1_94 delay_fixed_32_0_1_94_2984 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3002:142
    .clock (clock),
    .reset (reset),
    .in    (_dup279__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:425:111
    .out   (_delay_fixed_32_0_1_94_2984_out)
  );
  delay_fixed_32_0_1_70 delay_fixed_32_0_1_70_2985 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3003:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1019__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1165:116
    .out   (_delay_fixed_32_0_1_70_2985_out)
  );
  delay_fixed_32_0_1_1404 delay_fixed_32_0_1_1404_2986 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3004:150
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_2080),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_1404_2986_out)
  );
  delay_fixed_32_0_1_6 delay_fixed_32_0_1_6_2987 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3005:138
    .clock (clock),
    .reset (reset),
    .in    (_dup881__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1027:111
    .out   (_delay_fixed_32_0_1_6_2987_out)
  );
  delay_fixed_32_0_1_399 delay_fixed_32_0_1_399_2988 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3006:146
    .clock (clock),
    .reset (reset),
    .in    (_dup284__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:430:111
    .out   (_delay_fixed_32_0_1_399_2988_out)
  );
  delay_fixed_32_0_1_4 delay_fixed_32_0_1_4_2989 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3007:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1016__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1162:116
    .out   (_delay_fixed_32_0_1_4_2989_out)
  );
  delay_fixed_32_0_1_4 delay_fixed_32_0_1_4_2990 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3008:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1016__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1162:116
    .out   (_delay_fixed_32_0_1_4_2990_out)
  );
  delay_fixed_32_0_1_99 delay_fixed_32_0_1_99_2991 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3009:142
    .clock (clock),
    .reset (reset),
    .in    (_dup876__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1022:111
    .out   (_delay_fixed_32_0_1_99_2991_out)
  );
  delay_fixed_32_0_1_99 delay_fixed_32_0_1_99_2992 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3010:142
    .clock (clock),
    .reset (reset),
    .in    (_dup876__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1022:111
    .out   (_delay_fixed_32_0_1_99_2992_out)
  );
  delay_fixed_32_0_1_480 delay_fixed_32_0_1_480_2993 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3011:146
    .clock (clock),
    .reset (reset),
    .in    (_dup289__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:435:111
    .out   (_delay_fixed_32_0_1_480_2993_out)
  );
  delay_fixed_32_0_1_1032 delay_fixed_32_0_1_1032_2994 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3012:150
    .clock (clock),
    .reset (reset),
    .in    (_dup49_const_fix_32_0_1__0000000000000235_2320),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
    .out   (_delay_fixed_32_0_1_1032_2994_out)
  );
  delay_fixed_32_0_1_130 delay_fixed_32_0_1_130_2995 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3013:146
    .clock (clock),
    .reset (reset),
    .in    (_dup872__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1018:111
    .out   (_delay_fixed_32_0_1_130_2995_out)
  );
  delay_fixed_32_0_1_461 delay_fixed_32_0_1_461_2996 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3014:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1008__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1154:136
    .out   (_delay_fixed_32_0_1_461_2996_out)
  );
  delay_fixed_32_0_1_90 delay_fixed_32_0_1_90_2997 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3015:142
    .clock (clock),
    .reset (reset),
    .in    (_dup294__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:440:111
    .out   (_delay_fixed_32_0_1_90_2997_out)
  );
  delay_fixed_32_0_1_206 delay_fixed_32_0_1_206_2998 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3016:146
    .clock (clock),
    .reset (reset),
    .in    (_dup868__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1014:111
    .out   (_delay_fixed_32_0_1_206_2998_out)
  );
  delay_fixed_1_0_0_25 delay_fixed_1_0_0_25_2999 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3017:138
    .clock (clock),
    .reset (reset),
    .in    (_LT2004__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2150:139
    .out   (_delay_fixed_1_0_0_25_2999_out)
  );
  delay_fixed_32_0_1_1501 delay_fixed_32_0_1_1501_3000 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3018:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4813),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1501_3000_out)
  );
  delay_fixed_32_0_1_689 delay_fixed_32_0_1_689_3001 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3019:146
    .clock (clock),
    .reset (reset),
    .in    (_dup45_const_fix_32_0_1__0000000000000235_2320),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
    .out   (_delay_fixed_32_0_1_689_3001_out)
  );
  delay_fixed_32_0_1_206 delay_fixed_32_0_1_206_3002 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3020:146
    .clock (clock),
    .reset (reset),
    .in    (_dup868__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1014:111
    .out   (_delay_fixed_32_0_1_206_3002_out)
  );
  delay_fixed_32_0_1_1421 delay_fixed_32_0_1_1421_3003 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3021:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4809),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1421_3003_out)
  );
  delay_fixed_32_0_1_966 delay_fixed_32_0_1_966_3004 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3022:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_2388),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_966_3004_out)
  );
  delay_fixed_32_0_1_45 delay_fixed_32_0_1_45_3005 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3023:142
    .clock (clock),
    .reset (reset),
    .in    (_dup2001__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2147:154
    .out   (_delay_fixed_32_0_1_45_3005_out)
  );
  delay_fixed_32_0_1_1500 delay_fixed_32_0_1_1500_3006 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3024:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4813),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1500_3006_out)
  );
  delay_fixed_32_0_1_1037 delay_fixed_32_0_1_1037_3007 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3025:150
    .clock (clock),
    .reset (reset),
    .in    (_dup43_const_fix_32_0_1__0000000000000235_2320),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
    .out   (_delay_fixed_32_0_1_1037_3007_out)
  );
  delay_fixed_32_0_1_1455 delay_fixed_32_0_1_1455_3008 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3026:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4809),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1455_3008_out)
  );
  delay_fixed_32_0_1_287 delay_fixed_32_0_1_287_3009 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3027:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1004__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1150:116
    .out   (_delay_fixed_32_0_1_287_3009_out)
  );
  delay_fixed_32_0_1_225 delay_fixed_32_0_1_225_3010 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3028:146
    .clock (clock),
    .reset (reset),
    .in    (_dup864__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1010:111
    .out   (_delay_fixed_32_0_1_225_3010_out)
  );
  delay_fixed_32_0_1_480 delay_fixed_32_0_1_480_3011 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3029:146
    .clock (clock),
    .reset (reset),
    .in    (_dup289__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:435:111
    .out   (_delay_fixed_32_0_1_480_3011_out)
  );
  delay_fixed_32_0_1_225 delay_fixed_32_0_1_225_3012 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3030:146
    .clock (clock),
    .reset (reset),
    .in    (_dup864__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1010:111
    .out   (_delay_fixed_32_0_1_225_3012_out)
  );
  delay_fixed_32_0_1_39 delay_fixed_32_0_1_39_3013 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3031:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1936__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2082:116
    .out   (_delay_fixed_32_0_1_39_3013_out)
  );
  delay_fixed_32_0_1_25 delay_fixed_32_0_1_25_3014 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3032:142
    .clock (clock),
    .reset (reset),
    .in    (_dup999__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1145:111
    .out   (_delay_fixed_32_0_1_25_3014_out)
  );
  delay_fixed_32_0_1_25 delay_fixed_32_0_1_25_3015 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3033:142
    .clock (clock),
    .reset (reset),
    .in    (_dup999__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1145:111
    .out   (_delay_fixed_32_0_1_25_3015_out)
  );
  delay_fixed_32_0_1_9 delay_fixed_32_0_1_9_3016 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3034:138
    .clock (clock),
    .reset (reset),
    .in    (_MUX1995__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2141:169
    .out   (_delay_fixed_32_0_1_9_3016_out)
  );
  delay_fixed_32_0_1_1753 delay_fixed_32_0_1_1753_3017 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3035:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4791),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1753_3017_out)
  );
  delay_fixed_32_0_1_159 delay_fixed_32_0_1_159_3018 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3036:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL861__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1007:131
    .out   (_delay_fixed_32_0_1_159_3018_out)
  );
  delay_fixed_32_0_1_399 delay_fixed_32_0_1_399_3019 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3037:146
    .clock (clock),
    .reset (reset),
    .in    (_dup284__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:430:111
    .out   (_delay_fixed_32_0_1_399_3019_out)
  );
  delay_fixed_32_0_1_1677 delay_fixed_32_0_1_1677_3020 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3038:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4787),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1677_3020_out)
  );
  delay_fixed_32_0_1_757 delay_fixed_32_0_1_757_3021 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3039:146
    .clock (clock),
    .reset (reset),
    .in    (_dup49_const_fix_32_0_1__0000000000000235_1956),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
    .out   (_delay_fixed_32_0_1_757_3021_out)
  );
  delay_fixed_32_0_1_13 delay_fixed_32_0_1_13_3022 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3040:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1993__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2139:154
    .out   (_delay_fixed_32_0_1_13_3022_out)
  );
  delay_fixed_32_0_1_1724 delay_fixed_32_0_1_1724_3023 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3041:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4791),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1724_3023_out)
  );
  delay_fixed_32_0_1_1711 delay_fixed_32_0_1_1711_3024 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3042:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4787),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1711_3024_out)
  );
  delay_fixed_32_0_1_359 delay_fixed_32_0_1_359_3025 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3043:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL996__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1142:131
    .out   (_delay_fixed_32_0_1_359_3025_out)
  );
  delay_fixed_32_0_1_136 delay_fixed_32_0_1_136_3026 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3044:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL857__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1003:131
    .out   (_delay_fixed_32_0_1_136_3026_out)
  );
  delay_fixed_32_0_1_954 delay_fixed_32_0_1_954_3027 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3045:146
    .clock (clock),
    .reset (reset),
    .in    (_dup33_const_fix_32_0_1__0000000000000235_2320),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
    .out   (_delay_fixed_32_0_1_954_3027_out)
  );
  delay_fixed_32_0_1_787 delay_fixed_32_0_1_787_3028 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3046:146
    .clock (clock),
    .reset (reset),
    .in    (_dup45_const_fix_32_0_1__0000000000000235_1956),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
    .out   (_delay_fixed_32_0_1_787_3028_out)
  );
  delay_fixed_32_0_1_94 delay_fixed_32_0_1_94_3029 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3047:142
    .clock (clock),
    .reset (reset),
    .in    (_dup279__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:425:111
    .out   (_delay_fixed_32_0_1_94_3029_out)
  );
  delay_fixed_32_0_1_822 delay_fixed_32_0_1_822_3030 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3048:146
    .clock (clock),
    .reset (reset),
    .in    (_dup43_const_fix_32_0_1__0000000000000235_1956),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
    .out   (_delay_fixed_32_0_1_822_3030_out)
  );
  delay_fixed_1_0_0_94 delay_fixed_1_0_0_94_3031 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3049:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1988__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2134:139
    .out   (_delay_fixed_1_0_0_94_3031_out)
  );
  delay_fixed_32_0_1_1825 delay_fixed_32_0_1_1825_3032 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3050:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4769),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1825_3032_out)
  );
  delay_fixed_32_0_1_983 delay_fixed_32_0_1_983_3033 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3051:146
    .clock (clock),
    .reset (reset),
    .in    (_dup29_const_fix_32_0_1__0000000000000235_2320),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
    .out   (_delay_fixed_32_0_1_983_3033_out)
  );
  delay_fixed_32_0_1_86 delay_fixed_32_0_1_86_3034 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3052:142
    .clock (clock),
    .reset (reset),
    .in    (_dup852__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:998:111
    .out   (_delay_fixed_32_0_1_86_3034_out)
  );
  delay_fixed_32_0_1_1680 delay_fixed_32_0_1_1680_3035 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3053:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4765),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1680_3035_out)
  );
  delay_fixed_32_0_1_1076 delay_fixed_32_0_1_1076_3036 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3054:150
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_2352),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_1076_3036_out)
  );
  delay_fixed_32_0_1_778 delay_fixed_32_0_1_778_3037 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3055:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_689),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_778_3037_out)
  );
  delay_fixed_32_0_1_69 delay_fixed_32_0_1_69_3038 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3056:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1985__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2131:154
    .out   (_delay_fixed_32_0_1_69_3038_out)
  );
  delay_fixed_32_0_1_1783 delay_fixed_32_0_1_1783_3039 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3057:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4769),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1783_3039_out)
  );
  delay_fixed_32_0_1_1099 delay_fixed_32_0_1_1099_3040 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3058:150
    .clock (clock),
    .reset (reset),
    .in    (_dup27_const_fix_32_0_1__0000000000000235_2320),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
    .out   (_delay_fixed_32_0_1_1099_3040_out)
  );
  delay_fixed_32_0_1_634 delay_fixed_32_0_1_634_3041 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3059:146
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_685),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_634_3041_out)
  );
  delay_fixed_32_0_1_1714 delay_fixed_32_0_1_1714_3042 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3060:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4765),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1714_3042_out)
  );
  delay_fixed_32_0_1_87 delay_fixed_32_0_1_87_3043 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3061:142
    .clock (clock),
    .reset (reset),
    .in    (_dup988__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1134:111
    .out   (_delay_fixed_32_0_1_87_3043_out)
  );
  delay_fixed_32_0_1_126 delay_fixed_32_0_1_126_3044 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3062:146
    .clock (clock),
    .reset (reset),
    .in    (_dup849__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:995:111
    .out   (_delay_fixed_32_0_1_126_3044_out)
  );
  delay_fixed_32_0_1_31 delay_fixed_32_0_1_31_3045 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3063:142
    .clock (clock),
    .reset (reset),
    .in    (_dup270__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:416:111
    .out   (_delay_fixed_32_0_1_31_3045_out)
  );
  delay_fixed_32_0_1_126 delay_fixed_32_0_1_126_3046 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3064:146
    .clock (clock),
    .reset (reset),
    .in    (_dup849__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:995:111
    .out   (_delay_fixed_32_0_1_126_3046_out)
  );
  delay_fixed_32_0_1_717 delay_fixed_32_0_1_717_3047 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3065:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_677),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_717_3047_out)
  );
  delay_fixed_32_0_1_346 delay_fixed_32_0_1_346_3048 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3066:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1955__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2101:116
    .out   (_delay_fixed_32_0_1_346_3048_out)
  );
  delay_fixed_32_0_1_574 delay_fixed_32_0_1_574_3049 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3067:146
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_673),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_574_3049_out)
  );
  delay_fixed_32_0_1_386 delay_fixed_32_0_1_386_3050 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3068:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL984__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1130:131
    .out   (_delay_fixed_32_0_1_386_3050_out)
  );
  delay_fixed_32_0_1_31 delay_fixed_32_0_1_31_3051 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3069:142
    .clock (clock),
    .reset (reset),
    .in    (_dup270__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:416:111
    .out   (_delay_fixed_32_0_1_31_3051_out)
  );
  delay_fixed_32_0_1_26 delay_fixed_32_0_1_26_3052 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3070:142
    .clock (clock),
    .reset (reset),
    .in    (_MUX1979__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2125:169
    .out   (_delay_fixed_32_0_1_26_3052_out)
  );
  delay_fixed_32_0_1_1377 delay_fixed_32_0_1_1377_3053 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3071:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4747),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1377_3053_out)
  );
  delay_fixed_32_0_1_861 delay_fixed_32_0_1_861_3054 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3072:146
    .clock (clock),
    .reset (reset),
    .in    (_dup21_const_fix_32_0_1__0000000000000235_2320),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
    .out   (_delay_fixed_32_0_1_861_3054_out)
  );
  delay_fixed_32_0_1_218 delay_fixed_32_0_1_218_3055 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3073:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL845__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:991:131
    .out   (_delay_fixed_32_0_1_218_3055_out)
  );
  delay_fixed_32_0_1_1293 delay_fixed_32_0_1_1293_3056 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3074:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_4743),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1293_3056_out)
  );
  delay_fixed_32_0_1_835 delay_fixed_32_0_1_835_3057 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3075:146
    .clock (clock),
    .reset (reset),
    .in    (_dup33_const_fix_32_0_1__0000000000000235_1956),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
    .out   (_delay_fixed_32_0_1_835_3057_out)
  );
  delay_fixed_32_0_1_43 delay_fixed_32_0_1_43_3058 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3076:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1977__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2123:154
    .out   (_delay_fixed_32_0_1_43_3058_out)
  );
  delay_fixed_32_0_1_1370 delay_fixed_32_0_1_1370_3059 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3077:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4747),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1370_3059_out)
  );
  delay_fixed_32_0_1_125 delay_fixed_32_0_1_125_3060 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3078:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL980__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1126:131
    .out   (_delay_fixed_32_0_1_125_3060_out)
  );
  delay_fixed_32_0_1_51 delay_fixed_32_0_1_51_3061 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3079:142
    .clock (clock),
    .reset (reset),
    .in    (_dup266__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:412:111
    .out   (_delay_fixed_32_0_1_51_3061_out)
  );
  delay_fixed_32_0_1_1327 delay_fixed_32_0_1_1327_3062 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3080:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_4743),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1327_3062_out)
  );
  delay_fixed_32_0_1_209 delay_fixed_32_0_1_209_3063 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3081:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL841__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:987:131
    .out   (_delay_fixed_32_0_1_209_3063_out)
  );
  delay_fixed_32_0_1_51 delay_fixed_32_0_1_51_3064 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3082:142
    .clock (clock),
    .reset (reset),
    .in    (_dup266__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:412:111
    .out   (_delay_fixed_32_0_1_51_3064_out)
  );
  delay_fixed_32_0_1_1100 delay_fixed_32_0_1_1100_3065 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3083:150
    .clock (clock),
    .reset (reset),
    .in    (_dup17_const_fix_32_0_1__0000000000000235_2320),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
    .out   (_delay_fixed_32_0_1_1100_3065_out)
  );
  delay_fixed_32_0_1_1070 delay_fixed_32_0_1_1070_3066 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3084:150
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_2324),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_1070_3066_out)
  );
  delay_fixed_32_0_1_749 delay_fixed_32_0_1_749_3067 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3085:146
    .clock (clock),
    .reset (reset),
    .in    (_dup29_const_fix_32_0_1__0000000000000235_1956),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
    .out   (_delay_fixed_32_0_1_749_3067_out)
  );
  delay_fixed_1_0_0_60 delay_fixed_1_0_0_60_3068 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3086:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1094__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1240:139
    .out   (_delay_fixed_1_0_0_60_3068_out)
  );
  delay_fixed_32_0_1_2172 delay_fixed_32_0_1_2172_3069 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3087:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2585),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_2172_3069_out)
  );
  delay_fixed_32_0_1_47 delay_fixed_32_0_1_47_3070 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3088:142
    .clock (clock),
    .reset (reset),
    .in    (_dup262__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:408:111
    .out   (_delay_fixed_32_0_1_47_3070_out)
  );
  delay_fixed_32_0_1_2042 delay_fixed_32_0_1_2042_3071 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3089:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2581),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_2042_3071_out)
  );
  delay_fixed_32_0_1_47 delay_fixed_32_0_1_47_3072 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3090:142
    .clock (clock),
    .reset (reset),
    .in    (_dup262__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:408:111
    .out   (_delay_fixed_32_0_1_47_3072_out)
  );
  delay_fixed_32_0_1_63 delay_fixed_32_0_1_63_3073 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3091:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1091__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1237:154
    .out   (_delay_fixed_32_0_1_63_3073_out)
  );
  delay_fixed_32_0_1_2139 delay_fixed_32_0_1_2139_3074 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3092:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2585),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_2139_3074_out)
  );
  delay_fixed_32_0_1_2076 delay_fixed_32_0_1_2076_3075 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3093:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2581),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_2076_3075_out)
  );
  delay_fixed_32_0_1_28 delay_fixed_32_0_1_28_3076 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3094:142
    .clock (clock),
    .reset (reset),
    .in    (_dup257__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:403:111
    .out   (_delay_fixed_32_0_1_28_3076_out)
  );
  delay_fixed_32_0_1_28 delay_fixed_32_0_1_28_3077 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3095:142
    .clock (clock),
    .reset (reset),
    .in    (_dup257__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:403:111
    .out   (_delay_fixed_32_0_1_28_3077_out)
  );
  delay_fixed_32_0_1_365 delay_fixed_32_0_1_365_3078 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3096:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1061__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1207:116
    .out   (_delay_fixed_32_0_1_365_3078_out)
  );
  delay_fixed_32_0_1_37 delay_fixed_32_0_1_37_3079 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3097:142
    .clock (clock),
    .reset (reset),
    .in    (_dup253__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:399:111
    .out   (_delay_fixed_32_0_1_37_3079_out)
  );
  delay_fixed_32_0_1_37 delay_fixed_32_0_1_37_3080 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3098:142
    .clock (clock),
    .reset (reset),
    .in    (_dup253__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:399:111
    .out   (_delay_fixed_32_0_1_37_3080_out)
  );
  delay_fixed_32_0_1_216 delay_fixed_32_0_1_216_3081 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3099:146
    .clock (clock),
    .reset (reset),
    .in    (_dup389__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:535:111
    .out   (_delay_fixed_32_0_1_216_3081_out)
  );
  delay_fixed_32_0_1_33 delay_fixed_32_0_1_33_3082 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3100:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL251__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:397:131
    .out   (_delay_fixed_32_0_1_33_3082_out)
  );
  delay_fixed_32_0_1_17 delay_fixed_32_0_1_17_3083 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3101:142
    .clock (clock),
    .reset (reset),
    .in    (_dup394__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:540:111
    .out   (_delay_fixed_32_0_1_17_3083_out)
  );
  delay_fixed_32_0_1_110 delay_fixed_32_0_1_110_3084 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3102:146
    .clock (clock),
    .reset (reset),
    .in    (_dup49_const_fix_32_0_1__0000000000000235_570),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
    .out   (_delay_fixed_32_0_1_110_3084_out)
  );
  delay_fixed_32_0_1_110 delay_fixed_32_0_1_110_3085 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3103:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL248__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:394:131
    .out   (_delay_fixed_32_0_1_110_3085_out)
  );
  delay_fixed_32_0_1_17 delay_fixed_32_0_1_17_3086 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3104:142
    .clock (clock),
    .reset (reset),
    .in    (_dup394__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:540:111
    .out   (_delay_fixed_32_0_1_17_3086_out)
  );
  delay_fixed_32_0_1_39 delay_fixed_32_0_1_39_3087 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3105:142
    .clock (clock),
    .reset (reset),
    .in    (_dup45_const_fix_32_0_1__0000000000000235_570),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
    .out   (_delay_fixed_32_0_1_39_3087_out)
  );
  delay_fixed_32_0_1_83 delay_fixed_32_0_1_83_3088 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3106:142
    .clock (clock),
    .reset (reset),
    .in    (_dup43_const_fix_32_0_1__0000000000000235_570),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
    .out   (_delay_fixed_32_0_1_83_3088_out)
  );
  delay_fixed_32_0_1_15 delay_fixed_32_0_1_15_3089 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3107:142
    .clock (clock),
    .reset (reset),
    .in    (_dup245__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:391:111
    .out   (_delay_fixed_32_0_1_15_3089_out)
  );
  delay_fixed_32_0_1_216 delay_fixed_32_0_1_216_3090 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3108:146
    .clock (clock),
    .reset (reset),
    .in    (_dup389__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:535:111
    .out   (_delay_fixed_32_0_1_216_3090_out)
  );
  delay_fixed_32_0_1_53 delay_fixed_32_0_1_53_3091 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3109:142
    .clock (clock),
    .reset (reset),
    .in    (_dup240__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:386:111
    .out   (_delay_fixed_32_0_1_53_3091_out)
  );
  delay_fixed_32_0_1_53 delay_fixed_32_0_1_53_3092 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3110:142
    .clock (clock),
    .reset (reset),
    .in    (_dup240__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:386:111
    .out   (_delay_fixed_32_0_1_53_3092_out)
  );
  delay_fixed_32_0_1_143 delay_fixed_32_0_1_143_3093 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3111:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL238__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:384:131
    .out   (_delay_fixed_32_0_1_143_3093_out)
  );
  delay_fixed_32_0_1_270 delay_fixed_32_0_1_270_3094 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3112:146
    .clock (clock),
    .reset (reset),
    .in    (_dup384__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:530:111
    .out   (_delay_fixed_32_0_1_270_3094_out)
  );
  delay_fixed_32_0_1_160 delay_fixed_32_0_1_160_3095 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3113:146
    .clock (clock),
    .reset (reset),
    .in    (_dup33_const_fix_32_0_1__0000000000000235_570),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
    .out   (_delay_fixed_32_0_1_160_3095_out)
  );
  delay_fixed_32_0_1_146 delay_fixed_32_0_1_146_3096 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3114:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL235__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:381:131
    .out   (_delay_fixed_32_0_1_146_3096_out)
  );
  delay_fixed_32_0_1_50 delay_fixed_32_0_1_50_3097 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3115:142
    .clock (clock),
    .reset (reset),
    .in    (_dup29_const_fix_32_0_1__0000000000000235_570),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
    .out   (_delay_fixed_32_0_1_50_3097_out)
  );
  delay_fixed_32_0_1_256 delay_fixed_32_0_1_256_3098 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3116:146
    .clock (clock),
    .reset (reset),
    .in    (_dup27_const_fix_32_0_1__0000000000000235_570),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
    .out   (_delay_fixed_32_0_1_256_3098_out)
  );
  delay_fixed_32_0_1_52 delay_fixed_32_0_1_52_3099 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3117:142
    .clock (clock),
    .reset (reset),
    .in    (_dup231__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:377:111
    .out   (_delay_fixed_32_0_1_52_3099_out)
  );
  delay_fixed_32_0_1_212 delay_fixed_32_0_1_212_3100 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3118:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL229__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:375:131
    .out   (_delay_fixed_32_0_1_212_3100_out)
  );
  delay_fixed_32_0_1_97 delay_fixed_32_0_1_97_3101 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3119:142
    .clock (clock),
    .reset (reset),
    .in    (_dup21_const_fix_32_0_1__0000000000000235_570),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
    .out   (_delay_fixed_32_0_1_97_3101_out)
  );
  delay_fixed_32_0_1_225 delay_fixed_32_0_1_225_3102 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3120:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL226__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:372:131
    .out   (_delay_fixed_32_0_1_225_3102_out)
  );
  delay_fixed_32_0_1_66 delay_fixed_32_0_1_66_3103 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3121:142
    .clock (clock),
    .reset (reset),
    .in    (_dup17_const_fix_32_0_1__0000000000000235_570),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
    .out   (_delay_fixed_32_0_1_66_3103_out)
  );
  delay_fixed_32_0_1_143 delay_fixed_32_0_1_143_3104 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3122:146
    .clock (clock),
    .reset (reset),
    .in    (_dup15_const_fix_32_0_1__0000000000000235_570),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
    .out   (_delay_fixed_32_0_1_143_3104_out)
  );
  delay_fixed_32_0_1_13 delay_fixed_32_0_1_13_3105 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3123:142
    .clock (clock),
    .reset (reset),
    .in    (_dup223__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:369:111
    .out   (_delay_fixed_32_0_1_13_3105_out)
  );
  delay_fixed_32_0_1_122 delay_fixed_32_0_1_122_3106 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3124:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1149__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1295:116
    .out   (_delay_fixed_32_0_1_122_3106_out)
  );
  delay_fixed_32_0_1_97 delay_fixed_32_0_1_97_3107 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3125:142
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_564),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_97_3107_out)
  );
  delay_fixed_32_0_1_31 delay_fixed_32_0_1_31_3108 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3126:142
    .clock (clock),
    .reset (reset),
    .in    (_dup179__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:325:111
    .out   (_delay_fixed_32_0_1_31_3108_out)
  );
  delay_fixed_32_0_1_461 delay_fixed_32_0_1_461_3109 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3127:146
    .clock (clock),
    .reset (reset),
    .in    (_dup184__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:330:111
    .out   (_delay_fixed_32_0_1_461_3109_out)
  );
  delay_fixed_32_0_1_184 delay_fixed_32_0_1_184_3110 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3128:146
    .clock (clock),
    .reset (reset),
    .in    (_dup189__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:335:111
    .out   (_delay_fixed_32_0_1_184_3110_out)
  );
  delay_fixed_32_0_1_110 delay_fixed_32_0_1_110_3111 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3129:146
    .clock (clock),
    .reset (reset),
    .in    (_dup195__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:341:111
    .out   (_delay_fixed_32_0_1_110_3111_out)
  );
  delay_fixed_32_0_1_110 delay_fixed_32_0_1_110_3112 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3130:146
    .clock (clock),
    .reset (reset),
    .in    (_dup195__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:341:111
    .out   (_delay_fixed_32_0_1_110_3112_out)
  );
  delay_fixed_32_0_1_184 delay_fixed_32_0_1_184_3113 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3131:146
    .clock (clock),
    .reset (reset),
    .in    (_dup189__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:335:111
    .out   (_delay_fixed_32_0_1_184_3113_out)
  );
  delay_fixed_32_0_1_461 delay_fixed_32_0_1_461_3114 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3132:146
    .clock (clock),
    .reset (reset),
    .in    (_dup184__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:330:111
    .out   (_delay_fixed_32_0_1_461_3114_out)
  );
  delay_fixed_32_0_1_31 delay_fixed_32_0_1_31_3115 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3133:142
    .clock (clock),
    .reset (reset),
    .in    (_dup179__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:325:111
    .out   (_delay_fixed_32_0_1_31_3115_out)
  );
  delay_fixed_32_0_1_624 delay_fixed_32_0_1_624_3116 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3134:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_458),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_624_3116_out)
  );
  delay_fixed_32_0_1_493 delay_fixed_32_0_1_493_3117 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3135:146
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_454),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_493_3117_out)
  );
  delay_fixed_32_0_1_124 delay_fixed_32_0_1_124_3118 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3136:146
    .clock (clock),
    .reset (reset),
    .in    (_dup170__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:316:111
    .out   (_delay_fixed_32_0_1_124_3118_out)
  );
  delay_fixed_32_0_1_636 delay_fixed_32_0_1_636_3119 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3137:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_446),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_636_3119_out)
  );
  delay_fixed_32_0_1_486 delay_fixed_32_0_1_486_3120 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3138:146
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_442),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_486_3120_out)
  );
  delay_fixed_32_0_1_124 delay_fixed_32_0_1_124_3121 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3139:146
    .clock (clock),
    .reset (reset),
    .in    (_dup170__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:316:111
    .out   (_delay_fixed_32_0_1_124_3121_out)
  );
  delay_fixed_32_0_1_14 delay_fixed_32_0_1_14_3122 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3140:142
    .clock (clock),
    .reset (reset),
    .in    (_dup165__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:311:111
    .out   (_delay_fixed_32_0_1_14_3122_out)
  );
  delay_fixed_32_0_1_14 delay_fixed_32_0_1_14_3123 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3141:142
    .clock (clock),
    .reset (reset),
    .in    (_dup165__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:311:111
    .out   (_delay_fixed_32_0_1_14_3123_out)
  );
  delay_fixed_32_0_1_41 delay_fixed_32_0_1_41_3124 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3142:142
    .clock (clock),
    .reset (reset),
    .in    (_dup162__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:308:111
    .out   (_delay_fixed_32_0_1_41_3124_out)
  );
  delay_fixed_32_0_1_41 delay_fixed_32_0_1_41_3125 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3143:142
    .clock (clock),
    .reset (reset),
    .in    (_dup162__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:308:111
    .out   (_delay_fixed_32_0_1_41_3125_out)
  );
  delay_fixed_32_0_1_24 delay_fixed_32_0_1_24_3126 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3144:142
    .clock (clock),
    .reset (reset),
    .in    (_dup157__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:303:111
    .out   (_delay_fixed_32_0_1_24_3126_out)
  );
  delay_fixed_32_0_1_24 delay_fixed_32_0_1_24_3127 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3145:142
    .clock (clock),
    .reset (reset),
    .in    (_dup157__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:303:111
    .out   (_delay_fixed_32_0_1_24_3127_out)
  );
  delay_fixed_32_0_1_51 delay_fixed_32_0_1_51_3128 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3146:142
    .clock (clock),
    .reset (reset),
    .in    (_dup153__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:299:111
    .out   (_delay_fixed_32_0_1_51_3128_out)
  );
  delay_fixed_32_0_1_51 delay_fixed_32_0_1_51_3129 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3147:142
    .clock (clock),
    .reset (reset),
    .in    (_dup153__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:299:111
    .out   (_delay_fixed_32_0_1_51_3129_out)
  );
  delay_fixed_32_0_1_98 delay_fixed_32_0_1_98_3130 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3148:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL151__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:297:131
    .out   (_delay_fixed_32_0_1_98_3130_out)
  );
  delay_fixed_32_0_1_156 delay_fixed_32_0_1_156_3131 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3149:146
    .clock (clock),
    .reset (reset),
    .in    (_dup49_const_fix_32_0_1__0000000000000235_339),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
    .out   (_delay_fixed_32_0_1_156_3131_out)
  );
  delay_fixed_32_0_1_172 delay_fixed_32_0_1_172_3132 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3150:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL148__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:294:131
    .out   (_delay_fixed_32_0_1_172_3132_out)
  );
  delay_fixed_32_0_1_9 delay_fixed_32_0_1_9_3133 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3151:138
    .clock (clock),
    .reset (reset),
    .in    (_dup45_const_fix_32_0_1__0000000000000235_339),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
    .out   (_delay_fixed_32_0_1_9_3133_out)
  );
  delay_fixed_32_0_1_190 delay_fixed_32_0_1_190_3134 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3152:146
    .clock (clock),
    .reset (reset),
    .in    (_dup43_const_fix_32_0_1__0000000000000235_339),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
    .out   (_delay_fixed_32_0_1_190_3134_out)
  );
  delay_fixed_32_0_1_91 delay_fixed_32_0_1_91_3135 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3153:142
    .clock (clock),
    .reset (reset),
    .in    (_dup145__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:291:111
    .out   (_delay_fixed_32_0_1_91_3135_out)
  );
  delay_fixed_32_0_1_162 delay_fixed_32_0_1_162_3136 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3154:146
    .clock (clock),
    .reset (reset),
    .in    (_dup141__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:287:111
    .out   (_delay_fixed_32_0_1_162_3136_out)
  );
  delay_fixed_32_0_1_162 delay_fixed_32_0_1_162_3137 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3155:146
    .clock (clock),
    .reset (reset),
    .in    (_dup141__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:287:111
    .out   (_delay_fixed_32_0_1_162_3137_out)
  );
  delay_fixed_32_0_1_138 delay_fixed_32_0_1_138_3138 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3156:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL138__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:284:131
    .out   (_delay_fixed_32_0_1_138_3138_out)
  );
  delay_fixed_32_0_1_62 delay_fixed_32_0_1_62_3139 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3157:142
    .clock (clock),
    .reset (reset),
    .in    (_dup33_const_fix_32_0_1__0000000000000235_339),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
    .out   (_delay_fixed_32_0_1_62_3139_out)
  );
  delay_fixed_32_0_1_98 delay_fixed_32_0_1_98_3140 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3158:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL135__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:281:131
    .out   (_delay_fixed_32_0_1_98_3140_out)
  );
  delay_fixed_32_0_1_26 delay_fixed_32_0_1_26_3141 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3159:142
    .clock (clock),
    .reset (reset),
    .in    (_dup29_const_fix_32_0_1__0000000000000235_339),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
    .out   (_delay_fixed_32_0_1_26_3141_out)
  );
  delay_fixed_32_0_1_178 delay_fixed_32_0_1_178_3142 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3160:146
    .clock (clock),
    .reset (reset),
    .in    (_dup27_const_fix_32_0_1__0000000000000235_339),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
    .out   (_delay_fixed_32_0_1_178_3142_out)
  );
  delay_fixed_32_0_1_22 delay_fixed_32_0_1_22_3143 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3161:142
    .clock (clock),
    .reset (reset),
    .in    (_dup132__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:278:111
    .out   (_delay_fixed_32_0_1_22_3143_out)
  );
  delay_fixed_32_0_1_27 delay_fixed_32_0_1_27_3144 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3162:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL129__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:275:131
    .out   (_delay_fixed_32_0_1_27_3144_out)
  );
  delay_fixed_32_0_1_107 delay_fixed_32_0_1_107_3145 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3163:146
    .clock (clock),
    .reset (reset),
    .in    (_dup21_const_fix_32_0_1__0000000000000235_339),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
    .out   (_delay_fixed_32_0_1_107_3145_out)
  );
  delay_fixed_1_0_0_30 delay_fixed_1_0_0_30_3146 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3164:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1086__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1232:139
    .out   (_delay_fixed_1_0_0_30_3146_out)
  );
  delay_fixed_32_0_1_1774 delay_fixed_32_0_1_1774_3147 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3165:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2563),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1774_3147_out)
  );
  delay_fixed_32_0_1_117 delay_fixed_32_0_1_117_3148 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3166:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL126__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:272:131
    .out   (_delay_fixed_32_0_1_117_3148_out)
  );
  delay_fixed_32_0_1_1679 delay_fixed_32_0_1_1679_3149 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3167:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2559),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1679_3149_out)
  );
  delay_fixed_32_0_1_71 delay_fixed_32_0_1_71_3150 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3168:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1083__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1229:154
    .out   (_delay_fixed_32_0_1_71_3150_out)
  );
  delay_fixed_32_0_1_1784 delay_fixed_32_0_1_1784_3151 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3169:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2563),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1784_3151_out)
  );
  delay_fixed_32_0_1_9 delay_fixed_32_0_1_9_3152 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3170:138
    .clock (clock),
    .reset (reset),
    .in    (_dup17_const_fix_32_0_1__0000000000000235_339),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
    .out   (_delay_fixed_32_0_1_9_3152_out)
  );
  delay_fixed_32_0_1_1713 delay_fixed_32_0_1_1713_3153 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3171:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2559),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1713_3153_out)
  );
  delay_fixed_32_0_1_73 delay_fixed_32_0_1_73_3154 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3172:142
    .clock (clock),
    .reset (reset),
    .in    (_dup15_const_fix_32_0_1__0000000000000235_339),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
    .out   (_delay_fixed_32_0_1_73_3154_out)
  );
  delay_fixed_32_0_1_54 delay_fixed_32_0_1_54_3155 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3173:142
    .clock (clock),
    .reset (reset),
    .in    (_dup122__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:268:111
    .out   (_delay_fixed_32_0_1_54_3155_out)
  );
  delay_fixed_32_0_1_156 delay_fixed_32_0_1_156_3156 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3174:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1071__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1217:116
    .out   (_delay_fixed_32_0_1_156_3156_out)
  );
  delay_fixed_32_0_1_113 delay_fixed_32_0_1_113_3157 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3175:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_333),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_113_3157_out)
  );
  delay_fixed_1_0_0_52 delay_fixed_1_0_0_52_3158 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3176:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1078__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1224:139
    .out   (_delay_fixed_1_0_0_52_3158_out)
  );
  delay_fixed_32_0_1_1895 delay_fixed_32_0_1_1895_3159 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3177:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2541),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1895_3159_out)
  );
  delay_fixed_32_0_1_1762 delay_fixed_32_0_1_1762_3160 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3178:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2537),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1762_3160_out)
  );
  delay_fixed_32_0_1_39 delay_fixed_32_0_1_39_3161 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3179:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1075__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1221:154
    .out   (_delay_fixed_32_0_1_39_3161_out)
  );
  delay_fixed_32_0_1_1835 delay_fixed_32_0_1_1835_3162 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3180:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2541),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1835_3162_out)
  );
  delay_fixed_32_0_1_1796 delay_fixed_32_0_1_1796_3163 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3181:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2537),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1796_3163_out)
  );
  delay_fixed_32_0_1_156 delay_fixed_32_0_1_156_3164 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3182:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1071__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1217:116
    .out   (_delay_fixed_32_0_1_156_3164_out)
  );
  delay_fixed_1_0_0_2 delay_fixed_1_0_0_2_3165 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3183:134
    .clock (clock),
    .reset (reset),
    .in    (_LT1068__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1214:139
    .out   (_delay_fixed_1_0_0_2_3165_out)
  );
  delay_fixed_32_0_1_2006 delay_fixed_32_0_1_2006_3166 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3184:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2519),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_2006_3166_out)
  );
  delay_fixed_32_0_1_1953 delay_fixed_32_0_1_1953_3167 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3185:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2515),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1953_3167_out)
  );
  delay_fixed_32_0_1_4 delay_fixed_32_0_1_4_3168 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3186:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1065__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1211:154
    .out   (_delay_fixed_32_0_1_4_3168_out)
  );
  delay_fixed_32_0_1_1991 delay_fixed_32_0_1_1991_3169 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3187:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2519),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1991_3169_out)
  );
  delay_fixed_32_0_1_46 delay_fixed_32_0_1_46_3170 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3188:142
    .clock (clock),
    .reset (reset),
    .in    (_dup79__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:225:106
    .out   (_delay_fixed_32_0_1_46_3170_out)
  );
  delay_fixed_32_0_1_1987 delay_fixed_32_0_1_1987_3171 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3189:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_2515),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1987_3171_out)
  );
  delay_fixed_32_0_1_232 delay_fixed_32_0_1_232_3172 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3190:146
    .clock (clock),
    .reset (reset),
    .in    (_dup84__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:230:106
    .out   (_delay_fixed_32_0_1_232_3172_out)
  );
  delay_fixed_32_0_1_365 delay_fixed_32_0_1_365_3173 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3191:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1061__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1207:116
    .out   (_delay_fixed_32_0_1_365_3173_out)
  );
  delay_fixed_32_0_1_139 delay_fixed_32_0_1_139_3174 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3192:146
    .clock (clock),
    .reset (reset),
    .in    (_dup89__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:235:106
    .out   (_delay_fixed_32_0_1_139_3174_out)
  );
  delay_fixed_1_0_0_85 delay_fixed_1_0_0_85_3175 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3193:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1058__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1204:139
    .out   (_delay_fixed_1_0_0_85_3175_out)
  );
  delay_fixed_32_0_1_2274 delay_fixed_32_0_1_2274_3176 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3194:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_2497),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_2274_3176_out)
  );
  delay_fixed_32_0_1_81 delay_fixed_32_0_1_81_3177 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3195:142
    .clock (clock),
    .reset (reset),
    .in    (_dup94__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:240:106
    .out   (_delay_fixed_32_0_1_81_3177_out)
  );
  delay_fixed_32_0_1_81 delay_fixed_32_0_1_81_3178 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3196:142
    .clock (clock),
    .reset (reset),
    .in    (_dup94__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:240:106
    .out   (_delay_fixed_32_0_1_81_3178_out)
  );
  delay_fixed_32_0_1_139 delay_fixed_32_0_1_139_3179 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3197:146
    .clock (clock),
    .reset (reset),
    .in    (_dup89__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:235:106
    .out   (_delay_fixed_32_0_1_139_3179_out)
  );
  delay_fixed_32_0_1_232 delay_fixed_32_0_1_232_3180 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3198:146
    .clock (clock),
    .reset (reset),
    .in    (_dup84__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:230:106
    .out   (_delay_fixed_32_0_1_232_3180_out)
  );
  delay_fixed_32_0_1_46 delay_fixed_32_0_1_46_3181 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3199:142
    .clock (clock),
    .reset (reset),
    .in    (_dup79__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:225:106
    .out   (_delay_fixed_32_0_1_46_3181_out)
  );
  delay_fixed_32_0_1_552 delay_fixed_32_0_1_552_3182 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3200:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_227),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_552_3182_out)
  );
  delay_fixed_32_0_1_461 delay_fixed_32_0_1_461_3183 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3201:146
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_223),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_461_3183_out)
  );
  delay_fixed_32_0_1_1 delay_fixed_32_0_1_1_3184 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3202:138
    .clock (clock),
    .reset (reset),
    .in    (_dup69__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:215:106
    .out   (_delay_fixed_32_0_1_1_3184_out)
  );
  delay_fixed_32_0_1_566 delay_fixed_32_0_1_566_3185 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3203:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_215),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_566_3185_out)
  );
  delay_fixed_32_0_1_484 delay_fixed_32_0_1_484_3186 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3204:146
    .clock (clock),
    .reset (reset),
    .in    (_dup71_const_fix_32_0_1__00000000000000b5_211),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:217:1606
    .out   (_delay_fixed_32_0_1_484_3186_out)
  );
  delay_fixed_32_0_1_1 delay_fixed_32_0_1_1_3187 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3205:138
    .clock (clock),
    .reset (reset),
    .in    (_dup69__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:215:106
    .out   (_delay_fixed_32_0_1_1_3187_out)
  );
  delay_fixed_32_0_1_205 delay_fixed_32_0_1_205_3188 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3206:146
    .clock (clock),
    .reset (reset),
    .in    (_dup64__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:210:106
    .out   (_delay_fixed_32_0_1_205_3188_out)
  );
  delay_fixed_32_0_1_205 delay_fixed_32_0_1_205_3189 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3207:146
    .clock (clock),
    .reset (reset),
    .in    (_dup64__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:210:106
    .out   (_delay_fixed_32_0_1_205_3189_out)
  );
  delay_fixed_32_0_1_178 delay_fixed_32_0_1_178_3190 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3208:146
    .clock (clock),
    .reset (reset),
    .in    (_dup60__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:206:106
    .out   (_delay_fixed_32_0_1_178_3190_out)
  );
  delay_fixed_32_0_1_178 delay_fixed_32_0_1_178_3191 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3209:146
    .clock (clock),
    .reset (reset),
    .in    (_dup60__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:206:106
    .out   (_delay_fixed_32_0_1_178_3191_out)
  );
  delay_fixed_32_0_1_22 delay_fixed_32_0_1_22_3192 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3210:142
    .clock (clock),
    .reset (reset),
    .in    (_dup56__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:202:106
    .out   (_delay_fixed_32_0_1_22_3192_out)
  );
  delay_fixed_32_0_1_19 delay_fixed_32_0_1_19_3193 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3211:142
    .clock (clock),
    .reset (reset),
    .in    (_MUX1514__dfc_wire_2108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1660:169
    .out   (_delay_fixed_32_0_1_19_3193_out)
  );
  delay_fixed_32_0_1_1774 delay_fixed_32_0_1_1774_3194 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3212:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3611),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1774_3194_out)
  );
  delay_fixed_32_0_1_22 delay_fixed_32_0_1_22_3195 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3213:142
    .clock (clock),
    .reset (reset),
    .in    (_dup56__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:202:106
    .out   (_delay_fixed_32_0_1_22_3195_out)
  );
  delay_fixed_32_0_1_1736 delay_fixed_32_0_1_1736_3196 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3214:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3607),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1736_3196_out)
  );
  delay_fixed_32_0_1_16 delay_fixed_32_0_1_16_3197 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3215:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1512__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1658:154
    .out   (_delay_fixed_32_0_1_16_3197_out)
  );
  delay_fixed_32_0_1_1786 delay_fixed_32_0_1_1786_3198 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3216:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3611),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1786_3198_out)
  );
  delay_fixed_32_0_1_1770 delay_fixed_32_0_1_1770_3199 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3217:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3607),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1770_3199_out)
  );
  delay_fixed_32_0_1_11 delay_fixed_32_0_1_11_3200 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3218:142
    .clock (clock),
    .reset (reset),
    .in    (_dup52__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:198:106
    .out   (_delay_fixed_32_0_1_11_3200_out)
  );
  delay_fixed_32_0_1_11 delay_fixed_32_0_1_11_3201 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3219:142
    .clock (clock),
    .reset (reset),
    .in    (_dup52__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:198:106
    .out   (_delay_fixed_32_0_1_11_3201_out)
  );
  delay_fixed_32_0_1_259 delay_fixed_32_0_1_259_3202 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3220:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1145__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1291:136
    .out   (_delay_fixed_32_0_1_259_3202_out)
  );
  delay_fixed_32_0_1_905 delay_fixed_32_0_1_905_3203 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3221:146
    .clock (clock),
    .reset (reset),
    .in    (_dup33_const_fix_32_0_1__0000000000000235_2684),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:179:842
    .out   (_delay_fixed_32_0_1_905_3203_out)
  );
  delay_fixed_32_0_1_77 delay_fixed_32_0_1_77_3204 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3222:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL50__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:196:126
    .out   (_delay_fixed_32_0_1_77_3204_out)
  );
  delay_fixed_32_0_1_157 delay_fixed_32_0_1_157_3205 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3223:146
    .clock (clock),
    .reset (reset),
    .in    (_dup49_const_fix_32_0_1__0000000000000235_108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:195:842
    .out   (_delay_fixed_32_0_1_157_3205_out)
  );
  delay_fixed_32_0_1_222 delay_fixed_32_0_1_222_3206 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3224:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1141__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1287:136
    .out   (_delay_fixed_32_0_1_222_3206_out)
  );
  delay_fixed_32_0_1_85 delay_fixed_32_0_1_85_3207 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3225:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL46__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:192:126
    .out   (_delay_fixed_32_0_1_85_3207_out)
  );
  delay_fixed_32_0_1_100 delay_fixed_32_0_1_100_3208 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3226:146
    .clock (clock),
    .reset (reset),
    .in    (_dup45_const_fix_32_0_1__0000000000000235_108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:191:842
    .out   (_delay_fixed_32_0_1_100_3208_out)
  );
  delay_fixed_32_0_1_188 delay_fixed_32_0_1_188_3209 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3227:146
    .clock (clock),
    .reset (reset),
    .in    (_dup43_const_fix_32_0_1__0000000000000235_108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:189:842
    .out   (_delay_fixed_32_0_1_188_3209_out)
  );
  delay_fixed_32_0_1_128 delay_fixed_32_0_1_128_3210 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3228:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL1012__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1158:136
    .out   (_delay_fixed_32_0_1_128_3210_out)
  );
  delay_fixed_32_0_1_130 delay_fixed_32_0_1_130_3211 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3229:146
    .clock (clock),
    .reset (reset),
    .in    (_dup872__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1018:111
    .out   (_delay_fixed_32_0_1_130_3211_out)
  );
  delay_fixed_32_0_1_90 delay_fixed_32_0_1_90_3212 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3230:142
    .clock (clock),
    .reset (reset),
    .in    (_dup294__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:440:111
    .out   (_delay_fixed_32_0_1_90_3212_out)
  );
  delay_fixed_32_0_1_1 delay_fixed_32_0_1_1_3213 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3231:138
    .clock (clock),
    .reset (reset),
    .in    (_dup41__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:187:106
    .out   (_delay_fixed_32_0_1_1_3213_out)
  );
  delay_fixed_32_0_1_340 delay_fixed_32_0_1_340_3214 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3232:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1508__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1654:116
    .out   (_delay_fixed_32_0_1_340_3214_out)
  );
  delay_fixed_1_0_0_15 delay_fixed_1_0_0_15_3215 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3233:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1533__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1679:139
    .out   (_delay_fixed_1_0_0_15_3215_out)
  );
  delay_fixed_32_0_1_1439 delay_fixed_32_0_1_1439_3216 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3234:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3655),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1439_3216_out)
  );
  delay_fixed_32_0_1_5 delay_fixed_32_0_1_5_3217 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3235:138
    .clock (clock),
    .reset (reset),
    .in    (_dup37__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:183:106
    .out   (_delay_fixed_32_0_1_5_3217_out)
  );
  delay_fixed_32_0_1_1377 delay_fixed_32_0_1_1377_3218 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3236:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3651),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1377_3218_out)
  );
  delay_fixed_32_0_1_5 delay_fixed_32_0_1_5_3219 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3237:138
    .clock (clock),
    .reset (reset),
    .in    (_dup37__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:183:106
    .out   (_delay_fixed_32_0_1_5_3219_out)
  );
  delay_fixed_32_0_1_6 delay_fixed_32_0_1_6_3220 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3238:138
    .clock (clock),
    .reset (reset),
    .in    (_dup1530__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1676:154
    .out   (_delay_fixed_32_0_1_6_3220_out)
  );
  delay_fixed_32_0_1_1417 delay_fixed_32_0_1_1417_3221 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3239:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3655),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1417_3221_out)
  );
  delay_fixed_32_0_1_1411 delay_fixed_32_0_1_1411_3222 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3240:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3651),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1411_3222_out)
  );
  delay_fixed_32_0_1_280 delay_fixed_32_0_1_280_3223 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3241:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL34__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:180:126
    .out   (_delay_fixed_32_0_1_280_3223_out)
  );
  delay_fixed_32_0_1_10 delay_fixed_32_0_1_10_3224 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3242:142
    .clock (clock),
    .reset (reset),
    .in    (_dup25__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:171:106
    .out   (_delay_fixed_32_0_1_10_3224_out)
  );
  delay_fixed_32_0_1_23 delay_fixed_32_0_1_23_3225 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3243:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1518__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1664:116
    .out   (_delay_fixed_32_0_1_23_3225_out)
  );
  delay_fixed_32_0_1_148 delay_fixed_32_0_1_148_3226 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3244:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL30__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:176:126
    .out   (_delay_fixed_32_0_1_148_3226_out)
  );
  delay_fixed_32_0_1_72 delay_fixed_32_0_1_72_3227 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3245:142
    .clock (clock),
    .reset (reset),
    .in    (_dup29_const_fix_32_0_1__0000000000000235_108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:175:842
    .out   (_delay_fixed_32_0_1_72_3227_out)
  );
  delay_fixed_32_0_1_342 delay_fixed_32_0_1_342_3228 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3246:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1945__dfc_wire_68_113),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:2091:116
    .out   (_delay_fixed_32_0_1_342_3228_out)
  );
  delay_fixed_32_0_1_246 delay_fixed_32_0_1_246_3229 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3247:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL992__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1138:131
    .out   (_delay_fixed_32_0_1_246_3229_out)
  );
  delay_fixed_32_0_1_741 delay_fixed_32_0_1_741_3230 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3248:146
    .clock (clock),
    .reset (reset),
    .in    (_dup827_const_fix_32_0_1__0000000000000004_2024),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:973:1257
    .out   (_delay_fixed_32_0_1_741_3230_out)
  );
  delay_fixed_32_0_1_230 delay_fixed_32_0_1_230_3231 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3249:146
    .clock (clock),
    .reset (reset),
    .in    (_dup27_const_fix_32_0_1__0000000000000235_108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:173:842
    .out   (_delay_fixed_32_0_1_230_3231_out)
  );
  delay_fixed_32_0_1_340 delay_fixed_32_0_1_340_3232 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3250:146
    .clock (clock),
    .reset (reset),
    .in    (_dup1508__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1654:116
    .out   (_delay_fixed_32_0_1_340_3232_out)
  );
  delay_fixed_32_0_1_140 delay_fixed_32_0_1_140_3233 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3251:146
    .clock (clock),
    .reset (reset),
    .in    (_dup25__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:171:106
    .out   (_delay_fixed_32_0_1_140_3233_out)
  );
  delay_fixed_1_0_0_92 delay_fixed_1_0_0_92_3234 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3252:138
    .clock (clock),
    .reset (reset),
    .in    (_LT1505__dfc_wire_2112),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1651:139
    .out   (_delay_fixed_1_0_0_92_3234_out)
  );
  delay_fixed_32_0_1_1715 delay_fixed_32_0_1_1715_3235 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3253:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3589),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1715_3235_out)
  );
  delay_fixed_32_0_1_93 delay_fixed_32_0_1_93_3236 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3254:142
    .clock (clock),
    .reset (reset),
    .in    (_MUL22__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:168:126
    .out   (_delay_fixed_32_0_1_93_3236_out)
  );
  delay_fixed_32_0_1_1609 delay_fixed_32_0_1_1609_3237 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3255:150
    .clock (clock),
    .reset (reset),
    .in    (_dup898_const_fix_32_0_1__00000000000000ff_3585),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1044:6353
    .out   (_delay_fixed_32_0_1_1609_3237_out)
  );
  delay_fixed_32_0_1_90 delay_fixed_32_0_1_90_3238 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3256:142
    .clock (clock),
    .reset (reset),
    .in    (_dup21_const_fix_32_0_1__0000000000000235_108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:167:842
    .out   (_delay_fixed_32_0_1_90_3238_out)
  );
  delay_fixed_32_0_1_55 delay_fixed_32_0_1_55_3239 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3257:142
    .clock (clock),
    .reset (reset),
    .in    (_dup1502__dfc_wire_2103_2110),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1648:154
    .out   (_delay_fixed_32_0_1_55_3239_out)
  );
  delay_fixed_32_0_1_1698 delay_fixed_32_0_1_1698_3240 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3258:150
    .clock (clock),
    .reset (reset),
    .in    (_dup895_const_fix_32_0_1__00000000000000ff_3589),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:1041:6353
    .out   (_delay_fixed_32_0_1_1698_3240_out)
  );
  delay_fixed_32_0_1_167 delay_fixed_32_0_1_167_3241 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3259:146
    .clock (clock),
    .reset (reset),
    .in    (_MUL18__dfc_wire_107),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:164:126
    .out   (_delay_fixed_32_0_1_167_3241_out)
  );
  delay_fixed_32_0_1_34 delay_fixed_32_0_1_34_3242 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3260:142
    .clock (clock),
    .reset (reset),
    .in    (_dup17_const_fix_32_0_1__0000000000000235_108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:163:842
    .out   (_delay_fixed_32_0_1_34_3242_out)
  );
  delay_fixed_32_0_1_70 delay_fixed_32_0_1_70_3243 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3261:142
    .clock (clock),
    .reset (reset),
    .in    (_dup15_const_fix_32_0_1__0000000000000235_108),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:161:842
    .out   (_delay_fixed_32_0_1_70_3243_out)
  );
  delay_fixed_32_0_1_12 delay_fixed_32_0_1_12_3244 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3262:142
    .clock (clock),
    .reset (reset),
    .in    (_dup12__dfc_wire_68_105),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:158:106
    .out   (_delay_fixed_32_0_1_12_3244_out)
  );
  delay_fixed_32_0_1_119 delay_fixed_32_0_1_119_3245 (	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:3263:146
    .clock (clock),
    .reset (reset),
    .in    (_dup10_const_fix_32_0_1__0000000000000080_102),	// /home/nikita/Desktop/work/utopia/output/test/dfc/idct/idctFir.mlir:156:1986
    .out   (_delay_fixed_32_0_1_119_3245_out)
  );
endmodule

