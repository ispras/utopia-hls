// external module ADD_2x1

// external module MUL_2x1

// external module delay_fixed_16_0_1_12

// external module delay_fixed_16_0_1_22

// external module delay_fixed_16_0_1_66

// external module delay_fixed_16_0_1_8

// external module sink_1x0

// external module source_0x1

