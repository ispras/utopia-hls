module OUT(

    clock,
    reset,
    x);

input [15:0] x;
input clock;
input reset;
wire [15:0] x;
endmodule //OUT
