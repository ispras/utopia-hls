module W3_add_W5(

    clock,
    reset,
    value);

output [15:0] value;
input clock;
input reset;
wire [15:0] value;
assign value = (2408+1609);
endmodule //W3_add_W5
